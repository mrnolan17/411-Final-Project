module wallace_mul(
input [31:0] a, b,
input [1:0] mulop,
output logic [63:0] f
);

logic p [31:0][31:0];                // Partial product array

logic [991:0] s, c;                 // intermediate sum and cout

logic [63:0] curr_product, q, w;

logic [31:0] x, y;



integer i,j;

always_comb begin
q = {1'b0, c[533], c[676], c[773], c[772], c[839], c[838], c[837], c[836], c[882], c[881], c[880], c[879], c[878], c[877], c[913], c[912], c[911], c[910], c[909], c[908], c[907], c[906], c[905], c[929], c[928], c[927], c[926], c[925], c[924], c[923], c[922], c[921], c[920], c[919], c[918], c[917], c[916], c[915], c[914], s[914], c[888], c[887], c[886], c[885], c[884], c[883], s[883], c[843], c[842], c[841], c[840], s[840], c[775], c[774], s[774], c[677], s[677], c[534], s[534], s[320], s[0], p[0][1], p[0][0]};

w = {1'b0, p[31][31], s[533], s[676], s[773], s[772], s[839], s[838], s[837], s[836], s[882], s[881], s[880], s[879], s[878], s[877], s[913], s[912], s[911], s[910], s[909], s[908], s[907], s[906], s[905], s[929], s[928], s[927], s[926], s[925], s[924], s[923], s[922], s[921], s[920], s[919], s[918], s[917], s[916], s[915], s[378], s[889], s[888], s[887], s[886], s[885], s[884], s[348], s[844], s[843], s[842], s[841], s[21], s[776], s[775], s[11], s[678], p[6][0], s[535], p[4][0], p[3][0], p[2][0], p[1][0], 1'b0};


unique case(mulop)
2'b01 : begin
f = (a[31] ^ b[31]) ? (~curr_product + 64'b1) : curr_product;
x = a[31] ? (~a + 32'b1) : a;
y = b[31] ? (~b + 32'b1) : b;
end
2'b10 : begin
f = (a[31]) ? (~curr_product + 64'b1) : curr_product;
x = a[31] ? (~a + 32'b1) : a;
y = b;
end
2'b11 : begin
f = curr_product;
x = a;
y = b;
end
default : begin
f = (a[31] ^ b[31]) ? (~curr_product + 64'b1) : curr_product;
x = a[31] ? (~a + 32'b1) : a;
y = b[31] ? (~b + 32'b1) : b;
end
endcase
end

always@(x, y) begin
// PPartial products
for (i = 0; i <= 31; i = i + 1)

for (j = 0; j <= 31; j = j + 1)

p[j][i] <= x[j] & y[i];
 
end

carry_lookahead_adder64 cla(.A(q), .B(w), .Sum(curr_product));

HA ha_0_1 (.sum(s[0]), .cout(c[0]), .a(p[0][2]), .b(p[1][1]));
FA fa_0_2 (.sum(s[1]), .cout(c[1]), .a(p[0][3]), .b(p[1][2]), .c(p[2][1]));
FA fa_0_3 (.sum(s[2]), .cout(c[2]), .a(p[0][4]), .b(p[1][3]), .c(p[2][2]));
FA fa_0_4 (.sum(s[3]), .cout(c[3]), .a(p[0][5]), .b(p[1][4]), .c(p[2][3]));
FA fa_0_5 (.sum(s[4]), .cout(c[4]), .a(p[3][2]), .b(p[4][1]), .c(p[5][0]));
FA fa_0_6 (.sum(s[5]), .cout(c[5]), .a(p[0][6]), .b(p[1][5]), .c(p[2][4]));
FA fa_0_7 (.sum(s[6]), .cout(c[6]), .a(p[3][3]), .b(p[4][2]), .c(p[5][1]));
FA fa_0_8 (.sum(s[7]), .cout(c[7]), .a(p[0][7]), .b(p[1][6]), .c(p[2][5]));
FA fa_0_9 (.sum(s[8]), .cout(c[8]), .a(p[3][4]), .b(p[4][3]), .c(p[5][2]));
FA fa_0_10 (.sum(s[9]), .cout(c[9]), .a(p[0][8]), .b(p[1][7]), .c(p[2][6]));
FA fa_0_11 (.sum(s[10]), .cout(c[10]), .a(p[3][5]), .b(p[4][4]), .c(p[5][3]));
FA fa_0_12 (.sum(s[11]), .cout(c[11]), .a(p[6][2]), .b(p[7][1]), .c(p[8][0]));
FA fa_0_13 (.sum(s[12]), .cout(c[12]), .a(p[0][9]), .b(p[1][8]), .c(p[2][7]));
FA fa_0_14 (.sum(s[13]), .cout(c[13]), .a(p[3][6]), .b(p[4][5]), .c(p[5][4]));
FA fa_0_15 (.sum(s[14]), .cout(c[14]), .a(p[6][3]), .b(p[7][2]), .c(p[8][1]));
FA fa_0_16 (.sum(s[15]), .cout(c[15]), .a(p[0][10]), .b(p[1][9]), .c(p[2][8]));
FA fa_0_17 (.sum(s[16]), .cout(c[16]), .a(p[3][7]), .b(p[4][6]), .c(p[5][5]));
FA fa_0_18 (.sum(s[17]), .cout(c[17]), .a(p[6][4]), .b(p[7][3]), .c(p[8][2]));
FA fa_0_19 (.sum(s[18]), .cout(c[18]), .a(p[0][11]), .b(p[1][10]), .c(p[2][9]));
FA fa_0_20 (.sum(s[19]), .cout(c[19]), .a(p[3][8]), .b(p[4][7]), .c(p[5][6]));
FA fa_0_21 (.sum(s[20]), .cout(c[20]), .a(p[6][5]), .b(p[7][4]), .c(p[8][3]));
FA fa_0_22 (.sum(s[21]), .cout(c[21]), .a(p[9][2]), .b(p[10][1]), .c(p[11][0]));
FA fa_0_23 (.sum(s[22]), .cout(c[22]), .a(p[0][12]), .b(p[1][11]), .c(p[2][10]));
FA fa_0_24 (.sum(s[23]), .cout(c[23]), .a(p[3][9]), .b(p[4][8]), .c(p[5][7]));
FA fa_0_25 (.sum(s[24]), .cout(c[24]), .a(p[6][6]), .b(p[7][5]), .c(p[8][4]));
FA fa_0_26 (.sum(s[25]), .cout(c[25]), .a(p[9][3]), .b(p[10][2]), .c(p[11][1]));
FA fa_0_27 (.sum(s[26]), .cout(c[26]), .a(p[0][13]), .b(p[1][12]), .c(p[2][11]));
FA fa_0_28 (.sum(s[27]), .cout(c[27]), .a(p[3][10]), .b(p[4][9]), .c(p[5][8]));
FA fa_0_29 (.sum(s[28]), .cout(c[28]), .a(p[6][7]), .b(p[7][6]), .c(p[8][5]));
FA fa_0_30 (.sum(s[29]), .cout(c[29]), .a(p[9][4]), .b(p[10][3]), .c(p[11][2]));
FA fa_0_31 (.sum(s[30]), .cout(c[30]), .a(p[0][14]), .b(p[1][13]), .c(p[2][12]));
FA fa_0_32 (.sum(s[31]), .cout(c[31]), .a(p[3][11]), .b(p[4][10]), .c(p[5][9]));
FA fa_0_33 (.sum(s[32]), .cout(c[32]), .a(p[6][8]), .b(p[7][7]), .c(p[8][6]));
FA fa_0_34 (.sum(s[33]), .cout(c[33]), .a(p[9][5]), .b(p[10][4]), .c(p[11][3]));
FA fa_0_35 (.sum(s[34]), .cout(c[34]), .a(p[12][2]), .b(p[13][1]), .c(p[14][0]));
FA fa_0_36 (.sum(s[35]), .cout(c[35]), .a(p[0][15]), .b(p[1][14]), .c(p[2][13]));
FA fa_0_37 (.sum(s[36]), .cout(c[36]), .a(p[3][12]), .b(p[4][11]), .c(p[5][10]));
FA fa_0_38 (.sum(s[37]), .cout(c[37]), .a(p[6][9]), .b(p[7][8]), .c(p[8][7]));
FA fa_0_39 (.sum(s[38]), .cout(c[38]), .a(p[9][6]), .b(p[10][5]), .c(p[11][4]));
FA fa_0_40 (.sum(s[39]), .cout(c[39]), .a(p[12][3]), .b(p[13][2]), .c(p[14][1]));
FA fa_0_41 (.sum(s[40]), .cout(c[40]), .a(p[0][16]), .b(p[1][15]), .c(p[2][14]));
FA fa_0_42 (.sum(s[41]), .cout(c[41]), .a(p[3][13]), .b(p[4][12]), .c(p[5][11]));
FA fa_0_43 (.sum(s[42]), .cout(c[42]), .a(p[6][10]), .b(p[7][9]), .c(p[8][8]));
FA fa_0_44 (.sum(s[43]), .cout(c[43]), .a(p[9][7]), .b(p[10][6]), .c(p[11][5]));
FA fa_0_45 (.sum(s[44]), .cout(c[44]), .a(p[12][4]), .b(p[13][3]), .c(p[14][2]));
FA fa_0_46 (.sum(s[45]), .cout(c[45]), .a(p[0][17]), .b(p[1][16]), .c(p[2][15]));
FA fa_0_47 (.sum(s[46]), .cout(c[46]), .a(p[3][14]), .b(p[4][13]), .c(p[5][12]));
FA fa_0_48 (.sum(s[47]), .cout(c[47]), .a(p[6][11]), .b(p[7][10]), .c(p[8][9]));
FA fa_0_49 (.sum(s[48]), .cout(c[48]), .a(p[9][8]), .b(p[10][7]), .c(p[11][6]));
FA fa_0_50 (.sum(s[49]), .cout(c[49]), .a(p[12][5]), .b(p[13][4]), .c(p[14][3]));
FA fa_0_51 (.sum(s[50]), .cout(c[50]), .a(p[15][2]), .b(p[16][1]), .c(p[17][0]));
FA fa_0_52 (.sum(s[51]), .cout(c[51]), .a(p[0][18]), .b(p[1][17]), .c(p[2][16]));
FA fa_0_53 (.sum(s[52]), .cout(c[52]), .a(p[3][15]), .b(p[4][14]), .c(p[5][13]));
FA fa_0_54 (.sum(s[53]), .cout(c[53]), .a(p[6][12]), .b(p[7][11]), .c(p[8][10]));
FA fa_0_55 (.sum(s[54]), .cout(c[54]), .a(p[9][9]), .b(p[10][8]), .c(p[11][7]));
FA fa_0_56 (.sum(s[55]), .cout(c[55]), .a(p[12][6]), .b(p[13][5]), .c(p[14][4]));
FA fa_0_57 (.sum(s[56]), .cout(c[56]), .a(p[15][3]), .b(p[16][2]), .c(p[17][1]));
FA fa_0_58 (.sum(s[57]), .cout(c[57]), .a(p[0][19]), .b(p[1][18]), .c(p[2][17]));
FA fa_0_59 (.sum(s[58]), .cout(c[58]), .a(p[3][16]), .b(p[4][15]), .c(p[5][14]));
FA fa_0_60 (.sum(s[59]), .cout(c[59]), .a(p[6][13]), .b(p[7][12]), .c(p[8][11]));
FA fa_0_61 (.sum(s[60]), .cout(c[60]), .a(p[9][10]), .b(p[10][9]), .c(p[11][8]));
FA fa_0_62 (.sum(s[61]), .cout(c[61]), .a(p[12][7]), .b(p[13][6]), .c(p[14][5]));
FA fa_0_63 (.sum(s[62]), .cout(c[62]), .a(p[15][4]), .b(p[16][3]), .c(p[17][2]));
FA fa_0_64 (.sum(s[63]), .cout(c[63]), .a(p[0][20]), .b(p[1][19]), .c(p[2][18]));
FA fa_0_65 (.sum(s[64]), .cout(c[64]), .a(p[3][17]), .b(p[4][16]), .c(p[5][15]));
FA fa_0_66 (.sum(s[65]), .cout(c[65]), .a(p[6][14]), .b(p[7][13]), .c(p[8][12]));
FA fa_0_67 (.sum(s[66]), .cout(c[66]), .a(p[9][11]), .b(p[10][10]), .c(p[11][9]));
FA fa_0_68 (.sum(s[67]), .cout(c[67]), .a(p[12][8]), .b(p[13][7]), .c(p[14][6]));
FA fa_0_69 (.sum(s[68]), .cout(c[68]), .a(p[15][5]), .b(p[16][4]), .c(p[17][3]));
FA fa_0_70 (.sum(s[69]), .cout(c[69]), .a(p[18][2]), .b(p[19][1]), .c(p[20][0]));
FA fa_0_71 (.sum(s[70]), .cout(c[70]), .a(p[0][21]), .b(p[1][20]), .c(p[2][19]));
FA fa_0_72 (.sum(s[71]), .cout(c[71]), .a(p[3][18]), .b(p[4][17]), .c(p[5][16]));
FA fa_0_73 (.sum(s[72]), .cout(c[72]), .a(p[6][15]), .b(p[7][14]), .c(p[8][13]));
FA fa_0_74 (.sum(s[73]), .cout(c[73]), .a(p[9][12]), .b(p[10][11]), .c(p[11][10]));
FA fa_0_75 (.sum(s[74]), .cout(c[74]), .a(p[12][9]), .b(p[13][8]), .c(p[14][7]));
FA fa_0_76 (.sum(s[75]), .cout(c[75]), .a(p[15][6]), .b(p[16][5]), .c(p[17][4]));
FA fa_0_77 (.sum(s[76]), .cout(c[76]), .a(p[18][3]), .b(p[19][2]), .c(p[20][1]));
FA fa_0_78 (.sum(s[77]), .cout(c[77]), .a(p[0][22]), .b(p[1][21]), .c(p[2][20]));
FA fa_0_79 (.sum(s[78]), .cout(c[78]), .a(p[3][19]), .b(p[4][18]), .c(p[5][17]));
FA fa_0_80 (.sum(s[79]), .cout(c[79]), .a(p[6][16]), .b(p[7][15]), .c(p[8][14]));
FA fa_0_81 (.sum(s[80]), .cout(c[80]), .a(p[9][13]), .b(p[10][12]), .c(p[11][11]));
FA fa_0_82 (.sum(s[81]), .cout(c[81]), .a(p[12][10]), .b(p[13][9]), .c(p[14][8]));
FA fa_0_83 (.sum(s[82]), .cout(c[82]), .a(p[15][7]), .b(p[16][6]), .c(p[17][5]));
FA fa_0_84 (.sum(s[83]), .cout(c[83]), .a(p[18][4]), .b(p[19][3]), .c(p[20][2]));
FA fa_0_85 (.sum(s[84]), .cout(c[84]), .a(p[0][23]), .b(p[1][22]), .c(p[2][21]));
FA fa_0_86 (.sum(s[85]), .cout(c[85]), .a(p[3][20]), .b(p[4][19]), .c(p[5][18]));
FA fa_0_87 (.sum(s[86]), .cout(c[86]), .a(p[6][17]), .b(p[7][16]), .c(p[8][15]));
FA fa_0_88 (.sum(s[87]), .cout(c[87]), .a(p[9][14]), .b(p[10][13]), .c(p[11][12]));
FA fa_0_89 (.sum(s[88]), .cout(c[88]), .a(p[12][11]), .b(p[13][10]), .c(p[14][9]));
FA fa_0_90 (.sum(s[89]), .cout(c[89]), .a(p[15][8]), .b(p[16][7]), .c(p[17][6]));
FA fa_0_91 (.sum(s[90]), .cout(c[90]), .a(p[18][5]), .b(p[19][4]), .c(p[20][3]));
FA fa_0_92 (.sum(s[91]), .cout(c[91]), .a(p[21][2]), .b(p[22][1]), .c(p[23][0]));
FA fa_0_93 (.sum(s[92]), .cout(c[92]), .a(p[0][24]), .b(p[1][23]), .c(p[2][22]));
FA fa_0_94 (.sum(s[93]), .cout(c[93]), .a(p[3][21]), .b(p[4][20]), .c(p[5][19]));
FA fa_0_95 (.sum(s[94]), .cout(c[94]), .a(p[6][18]), .b(p[7][17]), .c(p[8][16]));
FA fa_0_96 (.sum(s[95]), .cout(c[95]), .a(p[9][15]), .b(p[10][14]), .c(p[11][13]));
FA fa_0_97 (.sum(s[96]), .cout(c[96]), .a(p[12][12]), .b(p[13][11]), .c(p[14][10]));
FA fa_0_98 (.sum(s[97]), .cout(c[97]), .a(p[15][9]), .b(p[16][8]), .c(p[17][7]));
FA fa_0_99 (.sum(s[98]), .cout(c[98]), .a(p[18][6]), .b(p[19][5]), .c(p[20][4]));
FA fa_0_100 (.sum(s[99]), .cout(c[99]), .a(p[21][3]), .b(p[22][2]), .c(p[23][1]));
FA fa_0_101 (.sum(s[100]), .cout(c[100]), .a(p[0][25]), .b(p[1][24]), .c(p[2][23]));
FA fa_0_102 (.sum(s[101]), .cout(c[101]), .a(p[3][22]), .b(p[4][21]), .c(p[5][20]));
FA fa_0_103 (.sum(s[102]), .cout(c[102]), .a(p[6][19]), .b(p[7][18]), .c(p[8][17]));
FA fa_0_104 (.sum(s[103]), .cout(c[103]), .a(p[9][16]), .b(p[10][15]), .c(p[11][14]));
FA fa_0_105 (.sum(s[104]), .cout(c[104]), .a(p[12][13]), .b(p[13][12]), .c(p[14][11]));
FA fa_0_106 (.sum(s[105]), .cout(c[105]), .a(p[15][10]), .b(p[16][9]), .c(p[17][8]));
FA fa_0_107 (.sum(s[106]), .cout(c[106]), .a(p[18][7]), .b(p[19][6]), .c(p[20][5]));
FA fa_0_108 (.sum(s[107]), .cout(c[107]), .a(p[21][4]), .b(p[22][3]), .c(p[23][2]));
FA fa_0_109 (.sum(s[108]), .cout(c[108]), .a(p[0][26]), .b(p[1][25]), .c(p[2][24]));
FA fa_0_110 (.sum(s[109]), .cout(c[109]), .a(p[3][23]), .b(p[4][22]), .c(p[5][21]));
FA fa_0_111 (.sum(s[110]), .cout(c[110]), .a(p[6][20]), .b(p[7][19]), .c(p[8][18]));
FA fa_0_112 (.sum(s[111]), .cout(c[111]), .a(p[9][17]), .b(p[10][16]), .c(p[11][15]));
FA fa_0_113 (.sum(s[112]), .cout(c[112]), .a(p[12][14]), .b(p[13][13]), .c(p[14][12]));
FA fa_0_114 (.sum(s[113]), .cout(c[113]), .a(p[15][11]), .b(p[16][10]), .c(p[17][9]));
FA fa_0_115 (.sum(s[114]), .cout(c[114]), .a(p[18][8]), .b(p[19][7]), .c(p[20][6]));
FA fa_0_116 (.sum(s[115]), .cout(c[115]), .a(p[21][5]), .b(p[22][4]), .c(p[23][3]));
FA fa_0_117 (.sum(s[116]), .cout(c[116]), .a(p[24][2]), .b(p[25][1]), .c(p[26][0]));
FA fa_0_118 (.sum(s[117]), .cout(c[117]), .a(p[0][27]), .b(p[1][26]), .c(p[2][25]));
FA fa_0_119 (.sum(s[118]), .cout(c[118]), .a(p[3][24]), .b(p[4][23]), .c(p[5][22]));
FA fa_0_120 (.sum(s[119]), .cout(c[119]), .a(p[6][21]), .b(p[7][20]), .c(p[8][19]));
FA fa_0_121 (.sum(s[120]), .cout(c[120]), .a(p[9][18]), .b(p[10][17]), .c(p[11][16]));
FA fa_0_122 (.sum(s[121]), .cout(c[121]), .a(p[12][15]), .b(p[13][14]), .c(p[14][13]));
FA fa_0_123 (.sum(s[122]), .cout(c[122]), .a(p[15][12]), .b(p[16][11]), .c(p[17][10]));
FA fa_0_124 (.sum(s[123]), .cout(c[123]), .a(p[18][9]), .b(p[19][8]), .c(p[20][7]));
FA fa_0_125 (.sum(s[124]), .cout(c[124]), .a(p[21][6]), .b(p[22][5]), .c(p[23][4]));
FA fa_0_126 (.sum(s[125]), .cout(c[125]), .a(p[24][3]), .b(p[25][2]), .c(p[26][1]));
FA fa_0_127 (.sum(s[126]), .cout(c[126]), .a(p[0][28]), .b(p[1][27]), .c(p[2][26]));
FA fa_0_128 (.sum(s[127]), .cout(c[127]), .a(p[3][25]), .b(p[4][24]), .c(p[5][23]));
FA fa_0_129 (.sum(s[128]), .cout(c[128]), .a(p[6][22]), .b(p[7][21]), .c(p[8][20]));
FA fa_0_130 (.sum(s[129]), .cout(c[129]), .a(p[9][19]), .b(p[10][18]), .c(p[11][17]));
FA fa_0_131 (.sum(s[130]), .cout(c[130]), .a(p[12][16]), .b(p[13][15]), .c(p[14][14]));
FA fa_0_132 (.sum(s[131]), .cout(c[131]), .a(p[15][13]), .b(p[16][12]), .c(p[17][11]));
FA fa_0_133 (.sum(s[132]), .cout(c[132]), .a(p[18][10]), .b(p[19][9]), .c(p[20][8]));
FA fa_0_134 (.sum(s[133]), .cout(c[133]), .a(p[21][7]), .b(p[22][6]), .c(p[23][5]));
FA fa_0_135 (.sum(s[134]), .cout(c[134]), .a(p[24][4]), .b(p[25][3]), .c(p[26][2]));
FA fa_0_136 (.sum(s[135]), .cout(c[135]), .a(p[0][29]), .b(p[1][28]), .c(p[2][27]));
FA fa_0_137 (.sum(s[136]), .cout(c[136]), .a(p[3][26]), .b(p[4][25]), .c(p[5][24]));
FA fa_0_138 (.sum(s[137]), .cout(c[137]), .a(p[6][23]), .b(p[7][22]), .c(p[8][21]));
FA fa_0_139 (.sum(s[138]), .cout(c[138]), .a(p[9][20]), .b(p[10][19]), .c(p[11][18]));
FA fa_0_140 (.sum(s[139]), .cout(c[139]), .a(p[12][17]), .b(p[13][16]), .c(p[14][15]));
FA fa_0_141 (.sum(s[140]), .cout(c[140]), .a(p[15][14]), .b(p[16][13]), .c(p[17][12]));
FA fa_0_142 (.sum(s[141]), .cout(c[141]), .a(p[18][11]), .b(p[19][10]), .c(p[20][9]));
FA fa_0_143 (.sum(s[142]), .cout(c[142]), .a(p[21][8]), .b(p[22][7]), .c(p[23][6]));
FA fa_0_144 (.sum(s[143]), .cout(c[143]), .a(p[24][5]), .b(p[25][4]), .c(p[26][3]));
FA fa_0_145 (.sum(s[144]), .cout(c[144]), .a(p[27][2]), .b(p[28][1]), .c(p[29][0]));
FA fa_0_146 (.sum(s[145]), .cout(c[145]), .a(p[0][30]), .b(p[1][29]), .c(p[2][28]));
FA fa_0_147 (.sum(s[146]), .cout(c[146]), .a(p[3][27]), .b(p[4][26]), .c(p[5][25]));
FA fa_0_148 (.sum(s[147]), .cout(c[147]), .a(p[6][24]), .b(p[7][23]), .c(p[8][22]));
FA fa_0_149 (.sum(s[148]), .cout(c[148]), .a(p[9][21]), .b(p[10][20]), .c(p[11][19]));
FA fa_0_150 (.sum(s[149]), .cout(c[149]), .a(p[12][18]), .b(p[13][17]), .c(p[14][16]));
FA fa_0_151 (.sum(s[150]), .cout(c[150]), .a(p[15][15]), .b(p[16][14]), .c(p[17][13]));
FA fa_0_152 (.sum(s[151]), .cout(c[151]), .a(p[18][12]), .b(p[19][11]), .c(p[20][10]));
FA fa_0_153 (.sum(s[152]), .cout(c[152]), .a(p[21][9]), .b(p[22][8]), .c(p[23][7]));
FA fa_0_154 (.sum(s[153]), .cout(c[153]), .a(p[24][6]), .b(p[25][5]), .c(p[26][4]));
FA fa_0_155 (.sum(s[154]), .cout(c[154]), .a(p[27][3]), .b(p[28][2]), .c(p[29][1]));
FA fa_0_156 (.sum(s[155]), .cout(c[155]), .a(p[0][31]), .b(p[1][30]), .c(p[2][29]));
FA fa_0_157 (.sum(s[156]), .cout(c[156]), .a(p[3][28]), .b(p[4][27]), .c(p[5][26]));
FA fa_0_158 (.sum(s[157]), .cout(c[157]), .a(p[6][25]), .b(p[7][24]), .c(p[8][23]));
FA fa_0_159 (.sum(s[158]), .cout(c[158]), .a(p[9][22]), .b(p[10][21]), .c(p[11][20]));
FA fa_0_160 (.sum(s[159]), .cout(c[159]), .a(p[12][19]), .b(p[13][18]), .c(p[14][17]));
FA fa_0_161 (.sum(s[160]), .cout(c[160]), .a(p[15][16]), .b(p[16][15]), .c(p[17][14]));
FA fa_0_162 (.sum(s[161]), .cout(c[161]), .a(p[18][13]), .b(p[19][12]), .c(p[20][11]));
FA fa_0_163 (.sum(s[162]), .cout(c[162]), .a(p[21][10]), .b(p[22][9]), .c(p[23][8]));
FA fa_0_164 (.sum(s[163]), .cout(c[163]), .a(p[24][7]), .b(p[25][6]), .c(p[26][5]));
FA fa_0_165 (.sum(s[164]), .cout(c[164]), .a(p[27][4]), .b(p[28][3]), .c(p[29][2]));
FA fa_0_166 (.sum(s[165]), .cout(c[165]), .a(p[1][31]), .b(p[2][30]), .c(p[3][29]));
FA fa_0_167 (.sum(s[166]), .cout(c[166]), .a(p[4][28]), .b(p[5][27]), .c(p[6][26]));
FA fa_0_168 (.sum(s[167]), .cout(c[167]), .a(p[7][25]), .b(p[8][24]), .c(p[9][23]));
FA fa_0_169 (.sum(s[168]), .cout(c[168]), .a(p[10][22]), .b(p[11][21]), .c(p[12][20]));
FA fa_0_170 (.sum(s[169]), .cout(c[169]), .a(p[13][19]), .b(p[14][18]), .c(p[15][17]));
FA fa_0_171 (.sum(s[170]), .cout(c[170]), .a(p[16][16]), .b(p[17][15]), .c(p[18][14]));
FA fa_0_172 (.sum(s[171]), .cout(c[171]), .a(p[19][13]), .b(p[20][12]), .c(p[21][11]));
FA fa_0_173 (.sum(s[172]), .cout(c[172]), .a(p[22][10]), .b(p[23][9]), .c(p[24][8]));
FA fa_0_174 (.sum(s[173]), .cout(c[173]), .a(p[25][7]), .b(p[26][6]), .c(p[27][5]));
FA fa_0_175 (.sum(s[174]), .cout(c[174]), .a(p[28][4]), .b(p[29][3]), .c(p[30][2]));
FA fa_0_176 (.sum(s[175]), .cout(c[175]), .a(p[2][31]), .b(p[3][30]), .c(p[4][29]));
FA fa_0_177 (.sum(s[176]), .cout(c[176]), .a(p[5][28]), .b(p[6][27]), .c(p[7][26]));
FA fa_0_178 (.sum(s[177]), .cout(c[177]), .a(p[8][25]), .b(p[9][24]), .c(p[10][23]));
FA fa_0_179 (.sum(s[178]), .cout(c[178]), .a(p[11][22]), .b(p[12][21]), .c(p[13][20]));
FA fa_0_180 (.sum(s[179]), .cout(c[179]), .a(p[14][19]), .b(p[15][18]), .c(p[16][17]));
FA fa_0_181 (.sum(s[180]), .cout(c[180]), .a(p[17][16]), .b(p[18][15]), .c(p[19][14]));
FA fa_0_182 (.sum(s[181]), .cout(c[181]), .a(p[20][13]), .b(p[21][12]), .c(p[22][11]));
FA fa_0_183 (.sum(s[182]), .cout(c[182]), .a(p[23][10]), .b(p[24][9]), .c(p[25][8]));
FA fa_0_184 (.sum(s[183]), .cout(c[183]), .a(p[26][7]), .b(p[27][6]), .c(p[28][5]));
FA fa_0_185 (.sum(s[184]), .cout(c[184]), .a(p[29][4]), .b(p[30][3]), .c(p[31][2]));
FA fa_0_186 (.sum(s[185]), .cout(c[185]), .a(p[3][31]), .b(p[4][30]), .c(p[5][29]));
FA fa_0_187 (.sum(s[186]), .cout(c[186]), .a(p[6][28]), .b(p[7][27]), .c(p[8][26]));
FA fa_0_188 (.sum(s[187]), .cout(c[187]), .a(p[9][25]), .b(p[10][24]), .c(p[11][23]));
FA fa_0_189 (.sum(s[188]), .cout(c[188]), .a(p[12][22]), .b(p[13][21]), .c(p[14][20]));
FA fa_0_190 (.sum(s[189]), .cout(c[189]), .a(p[15][19]), .b(p[16][18]), .c(p[17][17]));
FA fa_0_191 (.sum(s[190]), .cout(c[190]), .a(p[18][16]), .b(p[19][15]), .c(p[20][14]));
FA fa_0_192 (.sum(s[191]), .cout(c[191]), .a(p[21][13]), .b(p[22][12]), .c(p[23][11]));
FA fa_0_193 (.sum(s[192]), .cout(c[192]), .a(p[24][10]), .b(p[25][9]), .c(p[26][8]));
FA fa_0_194 (.sum(s[193]), .cout(c[193]), .a(p[27][7]), .b(p[28][6]), .c(p[29][5]));
FA fa_0_195 (.sum(s[194]), .cout(c[194]), .a(p[4][31]), .b(p[5][30]), .c(p[6][29]));
FA fa_0_196 (.sum(s[195]), .cout(c[195]), .a(p[7][28]), .b(p[8][27]), .c(p[9][26]));
FA fa_0_197 (.sum(s[196]), .cout(c[196]), .a(p[10][25]), .b(p[11][24]), .c(p[12][23]));
FA fa_0_198 (.sum(s[197]), .cout(c[197]), .a(p[13][22]), .b(p[14][21]), .c(p[15][20]));
FA fa_0_199 (.sum(s[198]), .cout(c[198]), .a(p[16][19]), .b(p[17][18]), .c(p[18][17]));
FA fa_0_200 (.sum(s[199]), .cout(c[199]), .a(p[19][16]), .b(p[20][15]), .c(p[21][14]));
FA fa_0_201 (.sum(s[200]), .cout(c[200]), .a(p[22][13]), .b(p[23][12]), .c(p[24][11]));
FA fa_0_202 (.sum(s[201]), .cout(c[201]), .a(p[25][10]), .b(p[26][9]), .c(p[27][8]));
FA fa_0_203 (.sum(s[202]), .cout(c[202]), .a(p[28][7]), .b(p[29][6]), .c(p[30][5]));
FA fa_0_204 (.sum(s[203]), .cout(c[203]), .a(p[5][31]), .b(p[6][30]), .c(p[7][29]));
FA fa_0_205 (.sum(s[204]), .cout(c[204]), .a(p[8][28]), .b(p[9][27]), .c(p[10][26]));
FA fa_0_206 (.sum(s[205]), .cout(c[205]), .a(p[11][25]), .b(p[12][24]), .c(p[13][23]));
FA fa_0_207 (.sum(s[206]), .cout(c[206]), .a(p[14][22]), .b(p[15][21]), .c(p[16][20]));
FA fa_0_208 (.sum(s[207]), .cout(c[207]), .a(p[17][19]), .b(p[18][18]), .c(p[19][17]));
FA fa_0_209 (.sum(s[208]), .cout(c[208]), .a(p[20][16]), .b(p[21][15]), .c(p[22][14]));
FA fa_0_210 (.sum(s[209]), .cout(c[209]), .a(p[23][13]), .b(p[24][12]), .c(p[25][11]));
FA fa_0_211 (.sum(s[210]), .cout(c[210]), .a(p[26][10]), .b(p[27][9]), .c(p[28][8]));
FA fa_0_212 (.sum(s[211]), .cout(c[211]), .a(p[29][7]), .b(p[30][6]), .c(p[31][5]));
FA fa_0_213 (.sum(s[212]), .cout(c[212]), .a(p[6][31]), .b(p[7][30]), .c(p[8][29]));
FA fa_0_214 (.sum(s[213]), .cout(c[213]), .a(p[9][28]), .b(p[10][27]), .c(p[11][26]));
FA fa_0_215 (.sum(s[214]), .cout(c[214]), .a(p[12][25]), .b(p[13][24]), .c(p[14][23]));
FA fa_0_216 (.sum(s[215]), .cout(c[215]), .a(p[15][22]), .b(p[16][21]), .c(p[17][20]));
FA fa_0_217 (.sum(s[216]), .cout(c[216]), .a(p[18][19]), .b(p[19][18]), .c(p[20][17]));
FA fa_0_218 (.sum(s[217]), .cout(c[217]), .a(p[21][16]), .b(p[22][15]), .c(p[23][14]));
FA fa_0_219 (.sum(s[218]), .cout(c[218]), .a(p[24][13]), .b(p[25][12]), .c(p[26][11]));
FA fa_0_220 (.sum(s[219]), .cout(c[219]), .a(p[27][10]), .b(p[28][9]), .c(p[29][8]));
FA fa_0_221 (.sum(s[220]), .cout(c[220]), .a(p[7][31]), .b(p[8][30]), .c(p[9][29]));
FA fa_0_222 (.sum(s[221]), .cout(c[221]), .a(p[10][28]), .b(p[11][27]), .c(p[12][26]));
FA fa_0_223 (.sum(s[222]), .cout(c[222]), .a(p[13][25]), .b(p[14][24]), .c(p[15][23]));
FA fa_0_224 (.sum(s[223]), .cout(c[223]), .a(p[16][22]), .b(p[17][21]), .c(p[18][20]));
FA fa_0_225 (.sum(s[224]), .cout(c[224]), .a(p[19][19]), .b(p[20][18]), .c(p[21][17]));
FA fa_0_226 (.sum(s[225]), .cout(c[225]), .a(p[22][16]), .b(p[23][15]), .c(p[24][14]));
FA fa_0_227 (.sum(s[226]), .cout(c[226]), .a(p[25][13]), .b(p[26][12]), .c(p[27][11]));
FA fa_0_228 (.sum(s[227]), .cout(c[227]), .a(p[28][10]), .b(p[29][9]), .c(p[30][8]));
FA fa_0_229 (.sum(s[228]), .cout(c[228]), .a(p[8][31]), .b(p[9][30]), .c(p[10][29]));
FA fa_0_230 (.sum(s[229]), .cout(c[229]), .a(p[11][28]), .b(p[12][27]), .c(p[13][26]));
FA fa_0_231 (.sum(s[230]), .cout(c[230]), .a(p[14][25]), .b(p[15][24]), .c(p[16][23]));
FA fa_0_232 (.sum(s[231]), .cout(c[231]), .a(p[17][22]), .b(p[18][21]), .c(p[19][20]));
FA fa_0_233 (.sum(s[232]), .cout(c[232]), .a(p[20][19]), .b(p[21][18]), .c(p[22][17]));
FA fa_0_234 (.sum(s[233]), .cout(c[233]), .a(p[23][16]), .b(p[24][15]), .c(p[25][14]));
FA fa_0_235 (.sum(s[234]), .cout(c[234]), .a(p[26][13]), .b(p[27][12]), .c(p[28][11]));
FA fa_0_236 (.sum(s[235]), .cout(c[235]), .a(p[29][10]), .b(p[30][9]), .c(p[31][8]));
FA fa_0_237 (.sum(s[236]), .cout(c[236]), .a(p[9][31]), .b(p[10][30]), .c(p[11][29]));
FA fa_0_238 (.sum(s[237]), .cout(c[237]), .a(p[12][28]), .b(p[13][27]), .c(p[14][26]));
FA fa_0_239 (.sum(s[238]), .cout(c[238]), .a(p[15][25]), .b(p[16][24]), .c(p[17][23]));
FA fa_0_240 (.sum(s[239]), .cout(c[239]), .a(p[18][22]), .b(p[19][21]), .c(p[20][20]));
FA fa_0_241 (.sum(s[240]), .cout(c[240]), .a(p[21][19]), .b(p[22][18]), .c(p[23][17]));
FA fa_0_242 (.sum(s[241]), .cout(c[241]), .a(p[24][16]), .b(p[25][15]), .c(p[26][14]));
FA fa_0_243 (.sum(s[242]), .cout(c[242]), .a(p[27][13]), .b(p[28][12]), .c(p[29][11]));
FA fa_0_244 (.sum(s[243]), .cout(c[243]), .a(p[10][31]), .b(p[11][30]), .c(p[12][29]));
FA fa_0_245 (.sum(s[244]), .cout(c[244]), .a(p[13][28]), .b(p[14][27]), .c(p[15][26]));
FA fa_0_246 (.sum(s[245]), .cout(c[245]), .a(p[16][25]), .b(p[17][24]), .c(p[18][23]));
FA fa_0_247 (.sum(s[246]), .cout(c[246]), .a(p[19][22]), .b(p[20][21]), .c(p[21][20]));
FA fa_0_248 (.sum(s[247]), .cout(c[247]), .a(p[22][19]), .b(p[23][18]), .c(p[24][17]));
FA fa_0_249 (.sum(s[248]), .cout(c[248]), .a(p[25][16]), .b(p[26][15]), .c(p[27][14]));
FA fa_0_250 (.sum(s[249]), .cout(c[249]), .a(p[28][13]), .b(p[29][12]), .c(p[30][11]));
FA fa_0_251 (.sum(s[250]), .cout(c[250]), .a(p[11][31]), .b(p[12][30]), .c(p[13][29]));
FA fa_0_252 (.sum(s[251]), .cout(c[251]), .a(p[14][28]), .b(p[15][27]), .c(p[16][26]));
FA fa_0_253 (.sum(s[252]), .cout(c[252]), .a(p[17][25]), .b(p[18][24]), .c(p[19][23]));
FA fa_0_254 (.sum(s[253]), .cout(c[253]), .a(p[20][22]), .b(p[21][21]), .c(p[22][20]));
FA fa_0_255 (.sum(s[254]), .cout(c[254]), .a(p[23][19]), .b(p[24][18]), .c(p[25][17]));
FA fa_0_256 (.sum(s[255]), .cout(c[255]), .a(p[26][16]), .b(p[27][15]), .c(p[28][14]));
FA fa_0_257 (.sum(s[256]), .cout(c[256]), .a(p[29][13]), .b(p[30][12]), .c(p[31][11]));
FA fa_0_258 (.sum(s[257]), .cout(c[257]), .a(p[12][31]), .b(p[13][30]), .c(p[14][29]));
FA fa_0_259 (.sum(s[258]), .cout(c[258]), .a(p[15][28]), .b(p[16][27]), .c(p[17][26]));
FA fa_0_260 (.sum(s[259]), .cout(c[259]), .a(p[18][25]), .b(p[19][24]), .c(p[20][23]));
FA fa_0_261 (.sum(s[260]), .cout(c[260]), .a(p[21][22]), .b(p[22][21]), .c(p[23][20]));
FA fa_0_262 (.sum(s[261]), .cout(c[261]), .a(p[24][19]), .b(p[25][18]), .c(p[26][17]));
FA fa_0_263 (.sum(s[262]), .cout(c[262]), .a(p[27][16]), .b(p[28][15]), .c(p[29][14]));
FA fa_0_264 (.sum(s[263]), .cout(c[263]), .a(p[13][31]), .b(p[14][30]), .c(p[15][29]));
FA fa_0_265 (.sum(s[264]), .cout(c[264]), .a(p[16][28]), .b(p[17][27]), .c(p[18][26]));
FA fa_0_266 (.sum(s[265]), .cout(c[265]), .a(p[19][25]), .b(p[20][24]), .c(p[21][23]));
FA fa_0_267 (.sum(s[266]), .cout(c[266]), .a(p[22][22]), .b(p[23][21]), .c(p[24][20]));
FA fa_0_268 (.sum(s[267]), .cout(c[267]), .a(p[25][19]), .b(p[26][18]), .c(p[27][17]));
FA fa_0_269 (.sum(s[268]), .cout(c[268]), .a(p[28][16]), .b(p[29][15]), .c(p[30][14]));
FA fa_0_270 (.sum(s[269]), .cout(c[269]), .a(p[14][31]), .b(p[15][30]), .c(p[16][29]));
FA fa_0_271 (.sum(s[270]), .cout(c[270]), .a(p[17][28]), .b(p[18][27]), .c(p[19][26]));
FA fa_0_272 (.sum(s[271]), .cout(c[271]), .a(p[20][25]), .b(p[21][24]), .c(p[22][23]));
FA fa_0_273 (.sum(s[272]), .cout(c[272]), .a(p[23][22]), .b(p[24][21]), .c(p[25][20]));
FA fa_0_274 (.sum(s[273]), .cout(c[273]), .a(p[26][19]), .b(p[27][18]), .c(p[28][17]));
FA fa_0_275 (.sum(s[274]), .cout(c[274]), .a(p[29][16]), .b(p[30][15]), .c(p[31][14]));
FA fa_0_276 (.sum(s[275]), .cout(c[275]), .a(p[15][31]), .b(p[16][30]), .c(p[17][29]));
FA fa_0_277 (.sum(s[276]), .cout(c[276]), .a(p[18][28]), .b(p[19][27]), .c(p[20][26]));
FA fa_0_278 (.sum(s[277]), .cout(c[277]), .a(p[21][25]), .b(p[22][24]), .c(p[23][23]));
FA fa_0_279 (.sum(s[278]), .cout(c[278]), .a(p[24][22]), .b(p[25][21]), .c(p[26][20]));
FA fa_0_280 (.sum(s[279]), .cout(c[279]), .a(p[27][19]), .b(p[28][18]), .c(p[29][17]));
FA fa_0_281 (.sum(s[280]), .cout(c[280]), .a(p[16][31]), .b(p[17][30]), .c(p[18][29]));
FA fa_0_282 (.sum(s[281]), .cout(c[281]), .a(p[19][28]), .b(p[20][27]), .c(p[21][26]));
FA fa_0_283 (.sum(s[282]), .cout(c[282]), .a(p[22][25]), .b(p[23][24]), .c(p[24][23]));
FA fa_0_284 (.sum(s[283]), .cout(c[283]), .a(p[25][22]), .b(p[26][21]), .c(p[27][20]));
FA fa_0_285 (.sum(s[284]), .cout(c[284]), .a(p[28][19]), .b(p[29][18]), .c(p[30][17]));
FA fa_0_286 (.sum(s[285]), .cout(c[285]), .a(p[17][31]), .b(p[18][30]), .c(p[19][29]));
FA fa_0_287 (.sum(s[286]), .cout(c[286]), .a(p[20][28]), .b(p[21][27]), .c(p[22][26]));
FA fa_0_288 (.sum(s[287]), .cout(c[287]), .a(p[23][25]), .b(p[24][24]), .c(p[25][23]));
FA fa_0_289 (.sum(s[288]), .cout(c[288]), .a(p[26][22]), .b(p[27][21]), .c(p[28][20]));
FA fa_0_290 (.sum(s[289]), .cout(c[289]), .a(p[29][19]), .b(p[30][18]), .c(p[31][17]));
FA fa_0_291 (.sum(s[290]), .cout(c[290]), .a(p[18][31]), .b(p[19][30]), .c(p[20][29]));
FA fa_0_292 (.sum(s[291]), .cout(c[291]), .a(p[21][28]), .b(p[22][27]), .c(p[23][26]));
FA fa_0_293 (.sum(s[292]), .cout(c[292]), .a(p[24][25]), .b(p[25][24]), .c(p[26][23]));
FA fa_0_294 (.sum(s[293]), .cout(c[293]), .a(p[27][22]), .b(p[28][21]), .c(p[29][20]));
FA fa_0_295 (.sum(s[294]), .cout(c[294]), .a(p[19][31]), .b(p[20][30]), .c(p[21][29]));
FA fa_0_296 (.sum(s[295]), .cout(c[295]), .a(p[22][28]), .b(p[23][27]), .c(p[24][26]));
FA fa_0_297 (.sum(s[296]), .cout(c[296]), .a(p[25][25]), .b(p[26][24]), .c(p[27][23]));
FA fa_0_298 (.sum(s[297]), .cout(c[297]), .a(p[28][22]), .b(p[29][21]), .c(p[30][20]));
FA fa_0_299 (.sum(s[298]), .cout(c[298]), .a(p[20][31]), .b(p[21][30]), .c(p[22][29]));
FA fa_0_300 (.sum(s[299]), .cout(c[299]), .a(p[23][28]), .b(p[24][27]), .c(p[25][26]));
FA fa_0_301 (.sum(s[300]), .cout(c[300]), .a(p[26][25]), .b(p[27][24]), .c(p[28][23]));
FA fa_0_302 (.sum(s[301]), .cout(c[301]), .a(p[29][22]), .b(p[30][21]), .c(p[31][20]));
FA fa_0_303 (.sum(s[302]), .cout(c[302]), .a(p[21][31]), .b(p[22][30]), .c(p[23][29]));
FA fa_0_304 (.sum(s[303]), .cout(c[303]), .a(p[24][28]), .b(p[25][27]), .c(p[26][26]));
FA fa_0_305 (.sum(s[304]), .cout(c[304]), .a(p[27][25]), .b(p[28][24]), .c(p[29][23]));
FA fa_0_306 (.sum(s[305]), .cout(c[305]), .a(p[22][31]), .b(p[23][30]), .c(p[24][29]));
FA fa_0_307 (.sum(s[306]), .cout(c[306]), .a(p[25][28]), .b(p[26][27]), .c(p[27][26]));
FA fa_0_308 (.sum(s[307]), .cout(c[307]), .a(p[28][25]), .b(p[29][24]), .c(p[30][23]));
FA fa_0_309 (.sum(s[308]), .cout(c[308]), .a(p[23][31]), .b(p[24][30]), .c(p[25][29]));
FA fa_0_310 (.sum(s[309]), .cout(c[309]), .a(p[26][28]), .b(p[27][27]), .c(p[28][26]));
FA fa_0_311 (.sum(s[310]), .cout(c[310]), .a(p[29][25]), .b(p[30][24]), .c(p[31][23]));
FA fa_0_312 (.sum(s[311]), .cout(c[311]), .a(p[24][31]), .b(p[25][30]), .c(p[26][29]));
FA fa_0_313 (.sum(s[312]), .cout(c[312]), .a(p[27][28]), .b(p[28][27]), .c(p[29][26]));
FA fa_0_314 (.sum(s[313]), .cout(c[313]), .a(p[25][31]), .b(p[26][30]), .c(p[27][29]));
FA fa_0_315 (.sum(s[314]), .cout(c[314]), .a(p[28][28]), .b(p[29][27]), .c(p[30][26]));
FA fa_0_316 (.sum(s[315]), .cout(c[315]), .a(p[26][31]), .b(p[27][30]), .c(p[28][29]));
FA fa_0_317 (.sum(s[316]), .cout(c[316]), .a(p[29][28]), .b(p[30][27]), .c(p[31][26]));
FA fa_0_318 (.sum(s[317]), .cout(c[317]), .a(p[27][31]), .b(p[28][30]), .c(p[29][29]));
FA fa_0_319 (.sum(s[318]), .cout(c[318]), .a(p[28][31]), .b(p[29][30]), .c(p[30][29]));
FA fa_0_320 (.sum(s[319]), .cout(c[319]), .a(p[29][31]), .b(p[30][30]), .c(p[31][29]));
HA ha_1_1 (.sum(s[320]), .cout(c[320]), .a(c[0]), .b(s[1]));
FA fa_1_2 (.sum(s[321]), .cout(c[321]), .a(c[1]), .b(s[2]), .c(p[3][1]));
FA fa_1_3 (.sum(s[322]), .cout(c[322]), .a(c[2]), .b(s[3]), .c(s[4]));
FA fa_1_4 (.sum(s[323]), .cout(c[323]), .a(c[3]), .b(c[4]), .c(s[5]));
FA fa_1_5 (.sum(s[324]), .cout(c[324]), .a(c[5]), .b(c[6]), .c(s[7]));
FA fa_1_6 (.sum(s[325]), .cout(c[325]), .a(s[8]), .b(p[6][1]), .c(p[7][0]));
FA fa_1_7 (.sum(s[326]), .cout(c[326]), .a(c[7]), .b(c[8]), .c(s[9]));
FA fa_1_8 (.sum(s[327]), .cout(c[327]), .a(c[9]), .b(c[10]), .c(c[11]));
FA fa_1_9 (.sum(s[328]), .cout(c[328]), .a(s[12]), .b(s[13]), .c(s[14]));
FA fa_1_10 (.sum(s[329]), .cout(c[329]), .a(c[12]), .b(c[13]), .c(c[14]));
FA fa_1_11 (.sum(s[330]), .cout(c[330]), .a(s[15]), .b(s[16]), .c(s[17]));
FA fa_1_12 (.sum(s[331]), .cout(c[331]), .a(c[15]), .b(c[16]), .c(c[17]));
FA fa_1_13 (.sum(s[332]), .cout(c[332]), .a(s[18]), .b(s[19]), .c(s[20]));
FA fa_1_14 (.sum(s[333]), .cout(c[333]), .a(c[18]), .b(c[19]), .c(c[20]));
FA fa_1_15 (.sum(s[334]), .cout(c[334]), .a(c[21]), .b(s[22]), .c(s[23]));
FA fa_1_16 (.sum(s[335]), .cout(c[335]), .a(s[24]), .b(s[25]), .c(p[12][0]));
FA fa_1_17 (.sum(s[336]), .cout(c[336]), .a(c[22]), .b(c[23]), .c(c[24]));
FA fa_1_18 (.sum(s[337]), .cout(c[337]), .a(c[25]), .b(s[26]), .c(s[27]));
FA fa_1_19 (.sum(s[338]), .cout(c[338]), .a(s[28]), .b(s[29]), .c(p[12][1]));
FA fa_1_20 (.sum(s[339]), .cout(c[339]), .a(c[26]), .b(c[27]), .c(c[28]));
FA fa_1_21 (.sum(s[340]), .cout(c[340]), .a(c[29]), .b(s[30]), .c(s[31]));
FA fa_1_22 (.sum(s[341]), .cout(c[341]), .a(s[32]), .b(s[33]), .c(s[34]));
FA fa_1_23 (.sum(s[342]), .cout(c[342]), .a(c[30]), .b(c[31]), .c(c[32]));
FA fa_1_24 (.sum(s[343]), .cout(c[343]), .a(c[33]), .b(c[34]), .c(s[35]));
FA fa_1_25 (.sum(s[344]), .cout(c[344]), .a(s[36]), .b(s[37]), .c(s[38]));
FA fa_1_26 (.sum(s[345]), .cout(c[345]), .a(c[35]), .b(c[36]), .c(c[37]));
FA fa_1_27 (.sum(s[346]), .cout(c[346]), .a(c[38]), .b(c[39]), .c(s[40]));
FA fa_1_28 (.sum(s[347]), .cout(c[347]), .a(s[41]), .b(s[42]), .c(s[43]));
FA fa_1_29 (.sum(s[348]), .cout(c[348]), .a(s[44]), .b(p[15][1]), .c(p[16][0]));
FA fa_1_30 (.sum(s[349]), .cout(c[349]), .a(c[40]), .b(c[41]), .c(c[42]));
FA fa_1_31 (.sum(s[350]), .cout(c[350]), .a(c[43]), .b(c[44]), .c(s[45]));
FA fa_1_32 (.sum(s[351]), .cout(c[351]), .a(s[46]), .b(s[47]), .c(s[48]));
FA fa_1_33 (.sum(s[352]), .cout(c[352]), .a(c[45]), .b(c[46]), .c(c[47]));
FA fa_1_34 (.sum(s[353]), .cout(c[353]), .a(c[48]), .b(c[49]), .c(c[50]));
FA fa_1_35 (.sum(s[354]), .cout(c[354]), .a(s[51]), .b(s[52]), .c(s[53]));
FA fa_1_36 (.sum(s[355]), .cout(c[355]), .a(s[54]), .b(s[55]), .c(s[56]));
FA fa_1_37 (.sum(s[356]), .cout(c[356]), .a(c[51]), .b(c[52]), .c(c[53]));
FA fa_1_38 (.sum(s[357]), .cout(c[357]), .a(c[54]), .b(c[55]), .c(c[56]));
FA fa_1_39 (.sum(s[358]), .cout(c[358]), .a(s[57]), .b(s[58]), .c(s[59]));
FA fa_1_40 (.sum(s[359]), .cout(c[359]), .a(s[60]), .b(s[61]), .c(s[62]));
FA fa_1_41 (.sum(s[360]), .cout(c[360]), .a(c[57]), .b(c[58]), .c(c[59]));
FA fa_1_42 (.sum(s[361]), .cout(c[361]), .a(c[60]), .b(c[61]), .c(c[62]));
FA fa_1_43 (.sum(s[362]), .cout(c[362]), .a(s[63]), .b(s[64]), .c(s[65]));
FA fa_1_44 (.sum(s[363]), .cout(c[363]), .a(s[66]), .b(s[67]), .c(s[68]));
FA fa_1_45 (.sum(s[364]), .cout(c[364]), .a(c[63]), .b(c[64]), .c(c[65]));
FA fa_1_46 (.sum(s[365]), .cout(c[365]), .a(c[66]), .b(c[67]), .c(c[68]));
FA fa_1_47 (.sum(s[366]), .cout(c[366]), .a(c[69]), .b(s[70]), .c(s[71]));
FA fa_1_48 (.sum(s[367]), .cout(c[367]), .a(s[72]), .b(s[73]), .c(s[74]));
FA fa_1_49 (.sum(s[368]), .cout(c[368]), .a(s[75]), .b(s[76]), .c(p[21][0]));
FA fa_1_50 (.sum(s[369]), .cout(c[369]), .a(c[70]), .b(c[71]), .c(c[72]));
FA fa_1_51 (.sum(s[370]), .cout(c[370]), .a(c[73]), .b(c[74]), .c(c[75]));
FA fa_1_52 (.sum(s[371]), .cout(c[371]), .a(c[76]), .b(s[77]), .c(s[78]));
FA fa_1_53 (.sum(s[372]), .cout(c[372]), .a(s[79]), .b(s[80]), .c(s[81]));
FA fa_1_54 (.sum(s[373]), .cout(c[373]), .a(s[82]), .b(s[83]), .c(p[21][1]));
FA fa_1_55 (.sum(s[374]), .cout(c[374]), .a(c[77]), .b(c[78]), .c(c[79]));
FA fa_1_56 (.sum(s[375]), .cout(c[375]), .a(c[80]), .b(c[81]), .c(c[82]));
FA fa_1_57 (.sum(s[376]), .cout(c[376]), .a(c[83]), .b(s[84]), .c(s[85]));
FA fa_1_58 (.sum(s[377]), .cout(c[377]), .a(s[86]), .b(s[87]), .c(s[88]));
FA fa_1_59 (.sum(s[378]), .cout(c[378]), .a(s[89]), .b(s[90]), .c(s[91]));
FA fa_1_60 (.sum(s[379]), .cout(c[379]), .a(c[84]), .b(c[85]), .c(c[86]));
FA fa_1_61 (.sum(s[380]), .cout(c[380]), .a(c[87]), .b(c[88]), .c(c[89]));
FA fa_1_62 (.sum(s[381]), .cout(c[381]), .a(c[90]), .b(c[91]), .c(s[92]));
FA fa_1_63 (.sum(s[382]), .cout(c[382]), .a(s[93]), .b(s[94]), .c(s[95]));
FA fa_1_64 (.sum(s[383]), .cout(c[383]), .a(s[96]), .b(s[97]), .c(s[98]));
FA fa_1_65 (.sum(s[384]), .cout(c[384]), .a(c[92]), .b(c[93]), .c(c[94]));
FA fa_1_66 (.sum(s[385]), .cout(c[385]), .a(c[95]), .b(c[96]), .c(c[97]));
FA fa_1_67 (.sum(s[386]), .cout(c[386]), .a(c[98]), .b(c[99]), .c(s[100]));
FA fa_1_68 (.sum(s[387]), .cout(c[387]), .a(s[101]), .b(s[102]), .c(s[103]));
FA fa_1_69 (.sum(s[388]), .cout(c[388]), .a(s[104]), .b(s[105]), .c(s[106]));
FA fa_1_70 (.sum(s[389]), .cout(c[389]), .a(s[107]), .b(p[24][1]), .c(p[25][0]));
FA fa_1_71 (.sum(s[390]), .cout(c[390]), .a(c[100]), .b(c[101]), .c(c[102]));
FA fa_1_72 (.sum(s[391]), .cout(c[391]), .a(c[103]), .b(c[104]), .c(c[105]));
FA fa_1_73 (.sum(s[392]), .cout(c[392]), .a(c[106]), .b(c[107]), .c(s[108]));
FA fa_1_74 (.sum(s[393]), .cout(c[393]), .a(s[109]), .b(s[110]), .c(s[111]));
FA fa_1_75 (.sum(s[394]), .cout(c[394]), .a(s[112]), .b(s[113]), .c(s[114]));
FA fa_1_76 (.sum(s[395]), .cout(c[395]), .a(c[108]), .b(c[109]), .c(c[110]));
FA fa_1_77 (.sum(s[396]), .cout(c[396]), .a(c[111]), .b(c[112]), .c(c[113]));
FA fa_1_78 (.sum(s[397]), .cout(c[397]), .a(c[114]), .b(c[115]), .c(c[116]));
FA fa_1_79 (.sum(s[398]), .cout(c[398]), .a(s[117]), .b(s[118]), .c(s[119]));
FA fa_1_80 (.sum(s[399]), .cout(c[399]), .a(s[120]), .b(s[121]), .c(s[122]));
FA fa_1_81 (.sum(s[400]), .cout(c[400]), .a(s[123]), .b(s[124]), .c(s[125]));
FA fa_1_82 (.sum(s[401]), .cout(c[401]), .a(c[117]), .b(c[118]), .c(c[119]));
FA fa_1_83 (.sum(s[402]), .cout(c[402]), .a(c[120]), .b(c[121]), .c(c[122]));
FA fa_1_84 (.sum(s[403]), .cout(c[403]), .a(c[123]), .b(c[124]), .c(c[125]));
FA fa_1_85 (.sum(s[404]), .cout(c[404]), .a(s[126]), .b(s[127]), .c(s[128]));
FA fa_1_86 (.sum(s[405]), .cout(c[405]), .a(s[129]), .b(s[130]), .c(s[131]));
FA fa_1_87 (.sum(s[406]), .cout(c[406]), .a(s[132]), .b(s[133]), .c(s[134]));
FA fa_1_88 (.sum(s[407]), .cout(c[407]), .a(c[126]), .b(c[127]), .c(c[128]));
FA fa_1_89 (.sum(s[408]), .cout(c[408]), .a(c[129]), .b(c[130]), .c(c[131]));
FA fa_1_90 (.sum(s[409]), .cout(c[409]), .a(c[132]), .b(c[133]), .c(c[134]));
FA fa_1_91 (.sum(s[410]), .cout(c[410]), .a(s[135]), .b(s[136]), .c(s[137]));
FA fa_1_92 (.sum(s[411]), .cout(c[411]), .a(s[138]), .b(s[139]), .c(s[140]));
FA fa_1_93 (.sum(s[412]), .cout(c[412]), .a(s[141]), .b(s[142]), .c(s[143]));
FA fa_1_94 (.sum(s[413]), .cout(c[413]), .a(c[135]), .b(c[136]), .c(c[137]));
FA fa_1_95 (.sum(s[414]), .cout(c[414]), .a(c[138]), .b(c[139]), .c(c[140]));
FA fa_1_96 (.sum(s[415]), .cout(c[415]), .a(c[141]), .b(c[142]), .c(c[143]));
FA fa_1_97 (.sum(s[416]), .cout(c[416]), .a(c[144]), .b(s[145]), .c(s[146]));
FA fa_1_98 (.sum(s[417]), .cout(c[417]), .a(s[147]), .b(s[148]), .c(s[149]));
FA fa_1_99 (.sum(s[418]), .cout(c[418]), .a(s[150]), .b(s[151]), .c(s[152]));
FA fa_1_100 (.sum(s[419]), .cout(c[419]), .a(s[153]), .b(s[154]), .c(p[30][0]));
FA fa_1_101 (.sum(s[420]), .cout(c[420]), .a(c[145]), .b(c[146]), .c(c[147]));
FA fa_1_102 (.sum(s[421]), .cout(c[421]), .a(c[148]), .b(c[149]), .c(c[150]));
FA fa_1_103 (.sum(s[422]), .cout(c[422]), .a(c[151]), .b(c[152]), .c(c[153]));
FA fa_1_104 (.sum(s[423]), .cout(c[423]), .a(c[154]), .b(s[155]), .c(s[156]));
FA fa_1_105 (.sum(s[424]), .cout(c[424]), .a(s[157]), .b(s[158]), .c(s[159]));
FA fa_1_106 (.sum(s[425]), .cout(c[425]), .a(s[160]), .b(s[161]), .c(s[162]));
FA fa_1_107 (.sum(s[426]), .cout(c[426]), .a(s[163]), .b(s[164]), .c(p[30][1]));
FA fa_1_108 (.sum(s[427]), .cout(c[427]), .a(c[155]), .b(c[156]), .c(c[157]));
FA fa_1_109 (.sum(s[428]), .cout(c[428]), .a(c[158]), .b(c[159]), .c(c[160]));
FA fa_1_110 (.sum(s[429]), .cout(c[429]), .a(c[161]), .b(c[162]), .c(c[163]));
FA fa_1_111 (.sum(s[430]), .cout(c[430]), .a(c[164]), .b(s[165]), .c(s[166]));
FA fa_1_112 (.sum(s[431]), .cout(c[431]), .a(s[167]), .b(s[168]), .c(s[169]));
FA fa_1_113 (.sum(s[432]), .cout(c[432]), .a(s[170]), .b(s[171]), .c(s[172]));
FA fa_1_114 (.sum(s[433]), .cout(c[433]), .a(s[173]), .b(s[174]), .c(p[31][1]));
FA fa_1_115 (.sum(s[434]), .cout(c[434]), .a(c[165]), .b(c[166]), .c(c[167]));
FA fa_1_116 (.sum(s[435]), .cout(c[435]), .a(c[168]), .b(c[169]), .c(c[170]));
FA fa_1_117 (.sum(s[436]), .cout(c[436]), .a(c[171]), .b(c[172]), .c(c[173]));
FA fa_1_118 (.sum(s[437]), .cout(c[437]), .a(c[174]), .b(s[175]), .c(s[176]));
FA fa_1_119 (.sum(s[438]), .cout(c[438]), .a(s[177]), .b(s[178]), .c(s[179]));
FA fa_1_120 (.sum(s[439]), .cout(c[439]), .a(s[180]), .b(s[181]), .c(s[182]));
FA fa_1_121 (.sum(s[440]), .cout(c[440]), .a(c[175]), .b(c[176]), .c(c[177]));
FA fa_1_122 (.sum(s[441]), .cout(c[441]), .a(c[178]), .b(c[179]), .c(c[180]));
FA fa_1_123 (.sum(s[442]), .cout(c[442]), .a(c[181]), .b(c[182]), .c(c[183]));
FA fa_1_124 (.sum(s[443]), .cout(c[443]), .a(c[184]), .b(s[185]), .c(s[186]));
FA fa_1_125 (.sum(s[444]), .cout(c[444]), .a(s[187]), .b(s[188]), .c(s[189]));
FA fa_1_126 (.sum(s[445]), .cout(c[445]), .a(s[190]), .b(s[191]), .c(s[192]));
FA fa_1_127 (.sum(s[446]), .cout(c[446]), .a(s[193]), .b(p[30][4]), .c(p[31][3]));
FA fa_1_128 (.sum(s[447]), .cout(c[447]), .a(c[185]), .b(c[186]), .c(c[187]));
FA fa_1_129 (.sum(s[448]), .cout(c[448]), .a(c[188]), .b(c[189]), .c(c[190]));
FA fa_1_130 (.sum(s[449]), .cout(c[449]), .a(c[191]), .b(c[192]), .c(c[193]));
FA fa_1_131 (.sum(s[450]), .cout(c[450]), .a(s[194]), .b(s[195]), .c(s[196]));
FA fa_1_132 (.sum(s[451]), .cout(c[451]), .a(s[197]), .b(s[198]), .c(s[199]));
FA fa_1_133 (.sum(s[452]), .cout(c[452]), .a(s[200]), .b(s[201]), .c(s[202]));
FA fa_1_134 (.sum(s[453]), .cout(c[453]), .a(c[194]), .b(c[195]), .c(c[196]));
FA fa_1_135 (.sum(s[454]), .cout(c[454]), .a(c[197]), .b(c[198]), .c(c[199]));
FA fa_1_136 (.sum(s[455]), .cout(c[455]), .a(c[200]), .b(c[201]), .c(c[202]));
FA fa_1_137 (.sum(s[456]), .cout(c[456]), .a(s[203]), .b(s[204]), .c(s[205]));
FA fa_1_138 (.sum(s[457]), .cout(c[457]), .a(s[206]), .b(s[207]), .c(s[208]));
FA fa_1_139 (.sum(s[458]), .cout(c[458]), .a(s[209]), .b(s[210]), .c(s[211]));
FA fa_1_140 (.sum(s[459]), .cout(c[459]), .a(c[203]), .b(c[204]), .c(c[205]));
FA fa_1_141 (.sum(s[460]), .cout(c[460]), .a(c[206]), .b(c[207]), .c(c[208]));
FA fa_1_142 (.sum(s[461]), .cout(c[461]), .a(c[209]), .b(c[210]), .c(c[211]));
FA fa_1_143 (.sum(s[462]), .cout(c[462]), .a(s[212]), .b(s[213]), .c(s[214]));
FA fa_1_144 (.sum(s[463]), .cout(c[463]), .a(s[215]), .b(s[216]), .c(s[217]));
FA fa_1_145 (.sum(s[464]), .cout(c[464]), .a(s[218]), .b(s[219]), .c(p[30][7]));
FA fa_1_146 (.sum(s[465]), .cout(c[465]), .a(c[212]), .b(c[213]), .c(c[214]));
FA fa_1_147 (.sum(s[466]), .cout(c[466]), .a(c[215]), .b(c[216]), .c(c[217]));
FA fa_1_148 (.sum(s[467]), .cout(c[467]), .a(c[218]), .b(c[219]), .c(s[220]));
FA fa_1_149 (.sum(s[468]), .cout(c[468]), .a(s[221]), .b(s[222]), .c(s[223]));
FA fa_1_150 (.sum(s[469]), .cout(c[469]), .a(s[224]), .b(s[225]), .c(s[226]));
FA fa_1_151 (.sum(s[470]), .cout(c[470]), .a(c[220]), .b(c[221]), .c(c[222]));
FA fa_1_152 (.sum(s[471]), .cout(c[471]), .a(c[223]), .b(c[224]), .c(c[225]));
FA fa_1_153 (.sum(s[472]), .cout(c[472]), .a(c[226]), .b(c[227]), .c(s[228]));
FA fa_1_154 (.sum(s[473]), .cout(c[473]), .a(s[229]), .b(s[230]), .c(s[231]));
FA fa_1_155 (.sum(s[474]), .cout(c[474]), .a(s[232]), .b(s[233]), .c(s[234]));
FA fa_1_156 (.sum(s[475]), .cout(c[475]), .a(c[228]), .b(c[229]), .c(c[230]));
FA fa_1_157 (.sum(s[476]), .cout(c[476]), .a(c[231]), .b(c[232]), .c(c[233]));
FA fa_1_158 (.sum(s[477]), .cout(c[477]), .a(c[234]), .b(c[235]), .c(s[236]));
FA fa_1_159 (.sum(s[478]), .cout(c[478]), .a(s[237]), .b(s[238]), .c(s[239]));
FA fa_1_160 (.sum(s[479]), .cout(c[479]), .a(s[240]), .b(s[241]), .c(s[242]));
FA fa_1_161 (.sum(s[480]), .cout(c[480]), .a(c[236]), .b(c[237]), .c(c[238]));
FA fa_1_162 (.sum(s[481]), .cout(c[481]), .a(c[239]), .b(c[240]), .c(c[241]));
FA fa_1_163 (.sum(s[482]), .cout(c[482]), .a(c[242]), .b(s[243]), .c(s[244]));
FA fa_1_164 (.sum(s[483]), .cout(c[483]), .a(s[245]), .b(s[246]), .c(s[247]));
FA fa_1_165 (.sum(s[484]), .cout(c[484]), .a(s[248]), .b(s[249]), .c(p[31][10]));
FA fa_1_166 (.sum(s[485]), .cout(c[485]), .a(c[243]), .b(c[244]), .c(c[245]));
FA fa_1_167 (.sum(s[486]), .cout(c[486]), .a(c[246]), .b(c[247]), .c(c[248]));
FA fa_1_168 (.sum(s[487]), .cout(c[487]), .a(c[249]), .b(s[250]), .c(s[251]));
FA fa_1_169 (.sum(s[488]), .cout(c[488]), .a(s[252]), .b(s[253]), .c(s[254]));
FA fa_1_170 (.sum(s[489]), .cout(c[489]), .a(c[250]), .b(c[251]), .c(c[252]));
FA fa_1_171 (.sum(s[490]), .cout(c[490]), .a(c[253]), .b(c[254]), .c(c[255]));
FA fa_1_172 (.sum(s[491]), .cout(c[491]), .a(c[256]), .b(s[257]), .c(s[258]));
FA fa_1_173 (.sum(s[492]), .cout(c[492]), .a(s[259]), .b(s[260]), .c(s[261]));
FA fa_1_174 (.sum(s[493]), .cout(c[493]), .a(s[262]), .b(p[30][13]), .c(p[31][12]));
FA fa_1_175 (.sum(s[494]), .cout(c[494]), .a(c[257]), .b(c[258]), .c(c[259]));
FA fa_1_176 (.sum(s[495]), .cout(c[495]), .a(c[260]), .b(c[261]), .c(c[262]));
FA fa_1_177 (.sum(s[496]), .cout(c[496]), .a(s[263]), .b(s[264]), .c(s[265]));
FA fa_1_178 (.sum(s[497]), .cout(c[497]), .a(s[266]), .b(s[267]), .c(s[268]));
FA fa_1_179 (.sum(s[498]), .cout(c[498]), .a(c[263]), .b(c[264]), .c(c[265]));
FA fa_1_180 (.sum(s[499]), .cout(c[499]), .a(c[266]), .b(c[267]), .c(c[268]));
FA fa_1_181 (.sum(s[500]), .cout(c[500]), .a(s[269]), .b(s[270]), .c(s[271]));
FA fa_1_182 (.sum(s[501]), .cout(c[501]), .a(s[272]), .b(s[273]), .c(s[274]));
FA fa_1_183 (.sum(s[502]), .cout(c[502]), .a(c[269]), .b(c[270]), .c(c[271]));
FA fa_1_184 (.sum(s[503]), .cout(c[503]), .a(c[272]), .b(c[273]), .c(c[274]));
FA fa_1_185 (.sum(s[504]), .cout(c[504]), .a(s[275]), .b(s[276]), .c(s[277]));
FA fa_1_186 (.sum(s[505]), .cout(c[505]), .a(s[278]), .b(s[279]), .c(p[30][16]));
FA fa_1_187 (.sum(s[506]), .cout(c[506]), .a(c[275]), .b(c[276]), .c(c[277]));
FA fa_1_188 (.sum(s[507]), .cout(c[507]), .a(c[278]), .b(c[279]), .c(s[280]));
FA fa_1_189 (.sum(s[508]), .cout(c[508]), .a(s[281]), .b(s[282]), .c(s[283]));
FA fa_1_190 (.sum(s[509]), .cout(c[509]), .a(c[280]), .b(c[281]), .c(c[282]));
FA fa_1_191 (.sum(s[510]), .cout(c[510]), .a(c[283]), .b(c[284]), .c(s[285]));
FA fa_1_192 (.sum(s[511]), .cout(c[511]), .a(s[286]), .b(s[287]), .c(s[288]));
FA fa_1_193 (.sum(s[512]), .cout(c[512]), .a(c[285]), .b(c[286]), .c(c[287]));
FA fa_1_194 (.sum(s[513]), .cout(c[513]), .a(c[288]), .b(c[289]), .c(s[290]));
FA fa_1_195 (.sum(s[514]), .cout(c[514]), .a(s[291]), .b(s[292]), .c(s[293]));
FA fa_1_196 (.sum(s[515]), .cout(c[515]), .a(c[290]), .b(c[291]), .c(c[292]));
FA fa_1_197 (.sum(s[516]), .cout(c[516]), .a(c[293]), .b(s[294]), .c(s[295]));
FA fa_1_198 (.sum(s[517]), .cout(c[517]), .a(s[296]), .b(s[297]), .c(p[31][19]));
FA fa_1_199 (.sum(s[518]), .cout(c[518]), .a(c[294]), .b(c[295]), .c(c[296]));
FA fa_1_200 (.sum(s[519]), .cout(c[519]), .a(c[297]), .b(s[298]), .c(s[299]));
FA fa_1_201 (.sum(s[520]), .cout(c[520]), .a(c[298]), .b(c[299]), .c(c[300]));
FA fa_1_202 (.sum(s[521]), .cout(c[521]), .a(c[301]), .b(s[302]), .c(s[303]));
FA fa_1_203 (.sum(s[522]), .cout(c[522]), .a(s[304]), .b(p[30][22]), .c(p[31][21]));
FA fa_1_204 (.sum(s[523]), .cout(c[523]), .a(c[302]), .b(c[303]), .c(c[304]));
FA fa_1_205 (.sum(s[524]), .cout(c[524]), .a(s[305]), .b(s[306]), .c(s[307]));
FA fa_1_206 (.sum(s[525]), .cout(c[525]), .a(c[305]), .b(c[306]), .c(c[307]));
FA fa_1_207 (.sum(s[526]), .cout(c[526]), .a(s[308]), .b(s[309]), .c(s[310]));
FA fa_1_208 (.sum(s[527]), .cout(c[527]), .a(c[308]), .b(c[309]), .c(c[310]));
FA fa_1_209 (.sum(s[528]), .cout(c[528]), .a(s[311]), .b(s[312]), .c(p[30][25]));
FA fa_1_210 (.sum(s[529]), .cout(c[529]), .a(c[311]), .b(c[312]), .c(s[313]));
FA fa_1_211 (.sum(s[530]), .cout(c[530]), .a(c[313]), .b(c[314]), .c(s[315]));
FA fa_1_212 (.sum(s[531]), .cout(c[531]), .a(c[315]), .b(c[316]), .c(s[317]));
FA fa_1_213 (.sum(s[532]), .cout(c[532]), .a(c[317]), .b(s[318]), .c(p[31][28]));
FA fa_1_214 (.sum(s[533]), .cout(c[533]), .a(c[319]), .b(p[30][31]), .c(p[31][30]));
HA ha_2_1 (.sum(s[534]), .cout(c[534]), .a(c[320]), .b(s[321]));
HA ha_2_2 (.sum(s[535]), .cout(c[535]), .a(c[321]), .b(s[322]));
FA fa_2_3 (.sum(s[536]), .cout(c[536]), .a(c[322]), .b(s[323]), .c(s[6]));
FA fa_2_4 (.sum(s[537]), .cout(c[537]), .a(c[323]), .b(s[324]), .c(s[325]));
FA fa_2_5 (.sum(s[538]), .cout(c[538]), .a(c[324]), .b(c[325]), .c(s[326]));
FA fa_2_6 (.sum(s[539]), .cout(c[539]), .a(c[326]), .b(s[327]), .c(s[328]));
FA fa_2_7 (.sum(s[540]), .cout(c[540]), .a(c[327]), .b(c[328]), .c(s[329]));
FA fa_2_8 (.sum(s[541]), .cout(c[541]), .a(s[330]), .b(p[9][1]), .c(p[10][0]));
FA fa_2_9 (.sum(s[542]), .cout(c[542]), .a(c[329]), .b(c[330]), .c(s[331]));
FA fa_2_10 (.sum(s[543]), .cout(c[543]), .a(c[331]), .b(c[332]), .c(s[333]));
FA fa_2_11 (.sum(s[544]), .cout(c[544]), .a(c[333]), .b(c[334]), .c(c[335]));
FA fa_2_12 (.sum(s[545]), .cout(c[545]), .a(s[336]), .b(s[337]), .c(s[338]));
FA fa_2_13 (.sum(s[546]), .cout(c[546]), .a(c[336]), .b(c[337]), .c(c[338]));
FA fa_2_14 (.sum(s[547]), .cout(c[547]), .a(s[339]), .b(s[340]), .c(s[341]));
FA fa_2_15 (.sum(s[548]), .cout(c[548]), .a(c[339]), .b(c[340]), .c(c[341]));
FA fa_2_16 (.sum(s[549]), .cout(c[549]), .a(s[342]), .b(s[343]), .c(s[344]));
FA fa_2_17 (.sum(s[550]), .cout(c[550]), .a(c[342]), .b(c[343]), .c(c[344]));
FA fa_2_18 (.sum(s[551]), .cout(c[551]), .a(s[345]), .b(s[346]), .c(s[347]));
FA fa_2_19 (.sum(s[552]), .cout(c[552]), .a(c[345]), .b(c[346]), .c(c[347]));
FA fa_2_20 (.sum(s[553]), .cout(c[553]), .a(c[348]), .b(s[349]), .c(s[350]));
FA fa_2_21 (.sum(s[554]), .cout(c[554]), .a(s[351]), .b(s[49]), .c(s[50]));
FA fa_2_22 (.sum(s[555]), .cout(c[555]), .a(c[349]), .b(c[350]), .c(c[351]));
FA fa_2_23 (.sum(s[556]), .cout(c[556]), .a(s[352]), .b(s[353]), .c(s[354]));
FA fa_2_24 (.sum(s[557]), .cout(c[557]), .a(c[352]), .b(c[353]), .c(c[354]));
FA fa_2_25 (.sum(s[558]), .cout(c[558]), .a(c[355]), .b(s[356]), .c(s[357]));
FA fa_2_26 (.sum(s[559]), .cout(c[559]), .a(s[358]), .b(s[359]), .c(p[18][1]));
FA fa_2_27 (.sum(s[560]), .cout(c[560]), .a(c[356]), .b(c[357]), .c(c[358]));
FA fa_2_28 (.sum(s[561]), .cout(c[561]), .a(c[359]), .b(s[360]), .c(s[361]));
FA fa_2_29 (.sum(s[562]), .cout(c[562]), .a(s[362]), .b(s[363]), .c(s[69]));
FA fa_2_30 (.sum(s[563]), .cout(c[563]), .a(c[360]), .b(c[361]), .c(c[362]));
FA fa_2_31 (.sum(s[564]), .cout(c[564]), .a(c[363]), .b(s[364]), .c(s[365]));
FA fa_2_32 (.sum(s[565]), .cout(c[565]), .a(s[366]), .b(s[367]), .c(s[368]));
FA fa_2_33 (.sum(s[566]), .cout(c[566]), .a(c[364]), .b(c[365]), .c(c[366]));
FA fa_2_34 (.sum(s[567]), .cout(c[567]), .a(c[367]), .b(c[368]), .c(s[369]));
FA fa_2_35 (.sum(s[568]), .cout(c[568]), .a(s[370]), .b(s[371]), .c(s[372]));
FA fa_2_36 (.sum(s[569]), .cout(c[569]), .a(c[369]), .b(c[370]), .c(c[371]));
FA fa_2_37 (.sum(s[570]), .cout(c[570]), .a(c[372]), .b(c[373]), .c(s[374]));
FA fa_2_38 (.sum(s[571]), .cout(c[571]), .a(s[375]), .b(s[376]), .c(s[377]));
FA fa_2_39 (.sum(s[572]), .cout(c[572]), .a(c[374]), .b(c[375]), .c(c[376]));
FA fa_2_40 (.sum(s[573]), .cout(c[573]), .a(c[377]), .b(c[378]), .c(s[379]));
FA fa_2_41 (.sum(s[574]), .cout(c[574]), .a(s[380]), .b(s[381]), .c(s[382]));
FA fa_2_42 (.sum(s[575]), .cout(c[575]), .a(s[383]), .b(s[99]), .c(p[24][0]));
FA fa_2_43 (.sum(s[576]), .cout(c[576]), .a(c[379]), .b(c[380]), .c(c[381]));
FA fa_2_44 (.sum(s[577]), .cout(c[577]), .a(c[382]), .b(c[383]), .c(s[384]));
FA fa_2_45 (.sum(s[578]), .cout(c[578]), .a(s[385]), .b(s[386]), .c(s[387]));
FA fa_2_46 (.sum(s[579]), .cout(c[579]), .a(c[384]), .b(c[385]), .c(c[386]));
FA fa_2_47 (.sum(s[580]), .cout(c[580]), .a(c[387]), .b(c[388]), .c(c[389]));
FA fa_2_48 (.sum(s[581]), .cout(c[581]), .a(s[390]), .b(s[391]), .c(s[392]));
FA fa_2_49 (.sum(s[582]), .cout(c[582]), .a(s[393]), .b(s[394]), .c(s[115]));
FA fa_2_50 (.sum(s[583]), .cout(c[583]), .a(c[390]), .b(c[391]), .c(c[392]));
FA fa_2_51 (.sum(s[584]), .cout(c[584]), .a(c[393]), .b(c[394]), .c(s[395]));
FA fa_2_52 (.sum(s[585]), .cout(c[585]), .a(s[396]), .b(s[397]), .c(s[398]));
FA fa_2_53 (.sum(s[586]), .cout(c[586]), .a(s[399]), .b(s[400]), .c(p[27][0]));
FA fa_2_54 (.sum(s[587]), .cout(c[587]), .a(c[395]), .b(c[396]), .c(c[397]));
FA fa_2_55 (.sum(s[588]), .cout(c[588]), .a(c[398]), .b(c[399]), .c(c[400]));
FA fa_2_56 (.sum(s[589]), .cout(c[589]), .a(s[401]), .b(s[402]), .c(s[403]));
FA fa_2_57 (.sum(s[590]), .cout(c[590]), .a(s[404]), .b(s[405]), .c(s[406]));
FA fa_2_58 (.sum(s[591]), .cout(c[591]), .a(c[401]), .b(c[402]), .c(c[403]));
FA fa_2_59 (.sum(s[592]), .cout(c[592]), .a(c[404]), .b(c[405]), .c(c[406]));
FA fa_2_60 (.sum(s[593]), .cout(c[593]), .a(s[407]), .b(s[408]), .c(s[409]));
FA fa_2_61 (.sum(s[594]), .cout(c[594]), .a(s[410]), .b(s[411]), .c(s[412]));
FA fa_2_62 (.sum(s[595]), .cout(c[595]), .a(c[407]), .b(c[408]), .c(c[409]));
FA fa_2_63 (.sum(s[596]), .cout(c[596]), .a(c[410]), .b(c[411]), .c(c[412]));
FA fa_2_64 (.sum(s[597]), .cout(c[597]), .a(s[413]), .b(s[414]), .c(s[415]));
FA fa_2_65 (.sum(s[598]), .cout(c[598]), .a(s[416]), .b(s[417]), .c(s[418]));
FA fa_2_66 (.sum(s[599]), .cout(c[599]), .a(c[413]), .b(c[414]), .c(c[415]));
FA fa_2_67 (.sum(s[600]), .cout(c[600]), .a(c[416]), .b(c[417]), .c(c[418]));
FA fa_2_68 (.sum(s[601]), .cout(c[601]), .a(c[419]), .b(s[420]), .c(s[421]));
FA fa_2_69 (.sum(s[602]), .cout(c[602]), .a(s[422]), .b(s[423]), .c(s[424]));
FA fa_2_70 (.sum(s[603]), .cout(c[603]), .a(s[425]), .b(s[426]), .c(p[31][0]));
FA fa_2_71 (.sum(s[604]), .cout(c[604]), .a(c[420]), .b(c[421]), .c(c[422]));
FA fa_2_72 (.sum(s[605]), .cout(c[605]), .a(c[423]), .b(c[424]), .c(c[425]));
FA fa_2_73 (.sum(s[606]), .cout(c[606]), .a(c[426]), .b(s[427]), .c(s[428]));
FA fa_2_74 (.sum(s[607]), .cout(c[607]), .a(s[429]), .b(s[430]), .c(s[431]));
FA fa_2_75 (.sum(s[608]), .cout(c[608]), .a(c[427]), .b(c[428]), .c(c[429]));
FA fa_2_76 (.sum(s[609]), .cout(c[609]), .a(c[430]), .b(c[431]), .c(c[432]));
FA fa_2_77 (.sum(s[610]), .cout(c[610]), .a(c[433]), .b(s[434]), .c(s[435]));
FA fa_2_78 (.sum(s[611]), .cout(c[611]), .a(s[436]), .b(s[437]), .c(s[438]));
FA fa_2_79 (.sum(s[612]), .cout(c[612]), .a(s[439]), .b(s[183]), .c(s[184]));
FA fa_2_80 (.sum(s[613]), .cout(c[613]), .a(c[434]), .b(c[435]), .c(c[436]));
FA fa_2_81 (.sum(s[614]), .cout(c[614]), .a(c[437]), .b(c[438]), .c(c[439]));
FA fa_2_82 (.sum(s[615]), .cout(c[615]), .a(s[440]), .b(s[441]), .c(s[442]));
FA fa_2_83 (.sum(s[616]), .cout(c[616]), .a(s[443]), .b(s[444]), .c(s[445]));
FA fa_2_84 (.sum(s[617]), .cout(c[617]), .a(c[440]), .b(c[441]), .c(c[442]));
FA fa_2_85 (.sum(s[618]), .cout(c[618]), .a(c[443]), .b(c[444]), .c(c[445]));
FA fa_2_86 (.sum(s[619]), .cout(c[619]), .a(c[446]), .b(s[447]), .c(s[448]));
FA fa_2_87 (.sum(s[620]), .cout(c[620]), .a(s[449]), .b(s[450]), .c(s[451]));
FA fa_2_88 (.sum(s[621]), .cout(c[621]), .a(c[447]), .b(c[448]), .c(c[449]));
FA fa_2_89 (.sum(s[622]), .cout(c[622]), .a(c[450]), .b(c[451]), .c(c[452]));
FA fa_2_90 (.sum(s[623]), .cout(c[623]), .a(s[453]), .b(s[454]), .c(s[455]));
FA fa_2_91 (.sum(s[624]), .cout(c[624]), .a(s[456]), .b(s[457]), .c(s[458]));
FA fa_2_92 (.sum(s[625]), .cout(c[625]), .a(c[453]), .b(c[454]), .c(c[455]));
FA fa_2_93 (.sum(s[626]), .cout(c[626]), .a(c[456]), .b(c[457]), .c(c[458]));
FA fa_2_94 (.sum(s[627]), .cout(c[627]), .a(s[459]), .b(s[460]), .c(s[461]));
FA fa_2_95 (.sum(s[628]), .cout(c[628]), .a(s[462]), .b(s[463]), .c(s[464]));
FA fa_2_96 (.sum(s[629]), .cout(c[629]), .a(c[459]), .b(c[460]), .c(c[461]));
FA fa_2_97 (.sum(s[630]), .cout(c[630]), .a(c[462]), .b(c[463]), .c(c[464]));
FA fa_2_98 (.sum(s[631]), .cout(c[631]), .a(s[465]), .b(s[466]), .c(s[467]));
FA fa_2_99 (.sum(s[632]), .cout(c[632]), .a(s[468]), .b(s[469]), .c(s[227]));
FA fa_2_100 (.sum(s[633]), .cout(c[633]), .a(c[465]), .b(c[466]), .c(c[467]));
FA fa_2_101 (.sum(s[634]), .cout(c[634]), .a(c[468]), .b(c[469]), .c(s[470]));
FA fa_2_102 (.sum(s[635]), .cout(c[635]), .a(s[471]), .b(s[472]), .c(s[473]));
FA fa_2_103 (.sum(s[636]), .cout(c[636]), .a(c[470]), .b(c[471]), .c(c[472]));
FA fa_2_104 (.sum(s[637]), .cout(c[637]), .a(c[473]), .b(c[474]), .c(s[475]));
FA fa_2_105 (.sum(s[638]), .cout(c[638]), .a(s[476]), .b(s[477]), .c(s[478]));
FA fa_2_106 (.sum(s[639]), .cout(c[639]), .a(s[479]), .b(p[30][10]), .c(p[31][9]));
FA fa_2_107 (.sum(s[640]), .cout(c[640]), .a(c[475]), .b(c[476]), .c(c[477]));
FA fa_2_108 (.sum(s[641]), .cout(c[641]), .a(c[478]), .b(c[479]), .c(s[480]));
FA fa_2_109 (.sum(s[642]), .cout(c[642]), .a(s[481]), .b(s[482]), .c(s[483]));
FA fa_2_110 (.sum(s[643]), .cout(c[643]), .a(c[480]), .b(c[481]), .c(c[482]));
FA fa_2_111 (.sum(s[644]), .cout(c[644]), .a(c[483]), .b(c[484]), .c(s[485]));
FA fa_2_112 (.sum(s[645]), .cout(c[645]), .a(s[486]), .b(s[487]), .c(s[488]));
FA fa_2_113 (.sum(s[646]), .cout(c[646]), .a(c[485]), .b(c[486]), .c(c[487]));
FA fa_2_114 (.sum(s[647]), .cout(c[647]), .a(c[488]), .b(s[489]), .c(s[490]));
FA fa_2_115 (.sum(s[648]), .cout(c[648]), .a(s[491]), .b(s[492]), .c(s[493]));
FA fa_2_116 (.sum(s[649]), .cout(c[649]), .a(c[489]), .b(c[490]), .c(c[491]));
FA fa_2_117 (.sum(s[650]), .cout(c[650]), .a(c[492]), .b(c[493]), .c(s[494]));
FA fa_2_118 (.sum(s[651]), .cout(c[651]), .a(s[495]), .b(s[496]), .c(s[497]));
FA fa_2_119 (.sum(s[652]), .cout(c[652]), .a(c[494]), .b(c[495]), .c(c[496]));
FA fa_2_120 (.sum(s[653]), .cout(c[653]), .a(c[497]), .b(s[498]), .c(s[499]));
FA fa_2_121 (.sum(s[654]), .cout(c[654]), .a(c[498]), .b(c[499]), .c(c[500]));
FA fa_2_122 (.sum(s[655]), .cout(c[655]), .a(c[501]), .b(s[502]), .c(s[503]));
FA fa_2_123 (.sum(s[656]), .cout(c[656]), .a(s[504]), .b(s[505]), .c(p[31][15]));
FA fa_2_124 (.sum(s[657]), .cout(c[657]), .a(c[502]), .b(c[503]), .c(c[504]));
FA fa_2_125 (.sum(s[658]), .cout(c[658]), .a(c[505]), .b(s[506]), .c(s[507]));
FA fa_2_126 (.sum(s[659]), .cout(c[659]), .a(s[508]), .b(s[284]), .c(p[31][16]));
FA fa_2_127 (.sum(s[660]), .cout(c[660]), .a(c[506]), .b(c[507]), .c(c[508]));
FA fa_2_128 (.sum(s[661]), .cout(c[661]), .a(s[509]), .b(s[510]), .c(s[511]));
FA fa_2_129 (.sum(s[662]), .cout(c[662]), .a(c[509]), .b(c[510]), .c(c[511]));
FA fa_2_130 (.sum(s[663]), .cout(c[663]), .a(s[512]), .b(s[513]), .c(s[514]));
FA fa_2_131 (.sum(s[664]), .cout(c[664]), .a(c[512]), .b(c[513]), .c(c[514]));
FA fa_2_132 (.sum(s[665]), .cout(c[665]), .a(s[515]), .b(s[516]), .c(s[517]));
FA fa_2_133 (.sum(s[666]), .cout(c[666]), .a(c[515]), .b(c[516]), .c(c[517]));
FA fa_2_134 (.sum(s[667]), .cout(c[667]), .a(s[518]), .b(s[519]), .c(s[300]));
FA fa_2_135 (.sum(s[668]), .cout(c[668]), .a(c[518]), .b(c[519]), .c(s[520]));
FA fa_2_136 (.sum(s[669]), .cout(c[669]), .a(c[520]), .b(c[521]), .c(c[522]));
FA fa_2_137 (.sum(s[670]), .cout(c[670]), .a(s[523]), .b(s[524]), .c(p[31][22]));
FA fa_2_138 (.sum(s[671]), .cout(c[671]), .a(c[523]), .b(c[524]), .c(s[525]));
FA fa_2_139 (.sum(s[672]), .cout(c[672]), .a(c[525]), .b(c[526]), .c(s[527]));
FA fa_2_140 (.sum(s[673]), .cout(c[673]), .a(c[527]), .b(c[528]), .c(s[529]));
FA fa_2_141 (.sum(s[674]), .cout(c[674]), .a(c[529]), .b(s[530]), .c(s[316]));
FA fa_2_142 (.sum(s[675]), .cout(c[675]), .a(c[530]), .b(s[531]), .c(p[30][28]));
FA fa_2_143 (.sum(s[676]), .cout(c[676]), .a(c[532]), .b(c[318]), .c(s[319]));
HA ha_3_1 (.sum(s[677]), .cout(c[677]), .a(c[535]), .b(s[536]));
HA ha_3_2 (.sum(s[678]), .cout(c[678]), .a(c[536]), .b(s[537]));
FA fa_3_3 (.sum(s[679]), .cout(c[679]), .a(c[537]), .b(s[538]), .c(s[10]));
FA fa_3_4 (.sum(s[680]), .cout(c[680]), .a(c[538]), .b(s[539]), .c(p[9][0]));
FA fa_3_5 (.sum(s[681]), .cout(c[681]), .a(c[539]), .b(s[540]), .c(s[541]));
FA fa_3_6 (.sum(s[682]), .cout(c[682]), .a(c[540]), .b(c[541]), .c(s[542]));
FA fa_3_7 (.sum(s[683]), .cout(c[683]), .a(c[542]), .b(s[543]), .c(s[334]));
FA fa_3_8 (.sum(s[684]), .cout(c[684]), .a(c[543]), .b(s[544]), .c(s[545]));
FA fa_3_9 (.sum(s[685]), .cout(c[685]), .a(c[544]), .b(c[545]), .c(s[546]));
FA fa_3_10 (.sum(s[686]), .cout(c[686]), .a(c[546]), .b(c[547]), .c(s[548]));
FA fa_3_11 (.sum(s[687]), .cout(c[687]), .a(s[549]), .b(s[39]), .c(p[15][0]));
FA fa_3_12 (.sum(s[688]), .cout(c[688]), .a(c[548]), .b(c[549]), .c(s[550]));
FA fa_3_13 (.sum(s[689]), .cout(c[689]), .a(c[550]), .b(c[551]), .c(s[552]));
FA fa_3_14 (.sum(s[690]), .cout(c[690]), .a(c[552]), .b(c[553]), .c(c[554]));
FA fa_3_15 (.sum(s[691]), .cout(c[691]), .a(s[555]), .b(s[556]), .c(s[355]));
FA fa_3_16 (.sum(s[692]), .cout(c[692]), .a(c[555]), .b(c[556]), .c(s[557]));
FA fa_3_17 (.sum(s[693]), .cout(c[693]), .a(s[558]), .b(s[559]), .c(p[19][0]));
FA fa_3_18 (.sum(s[694]), .cout(c[694]), .a(c[557]), .b(c[558]), .c(c[559]));
FA fa_3_19 (.sum(s[695]), .cout(c[695]), .a(s[560]), .b(s[561]), .c(s[562]));
FA fa_3_20 (.sum(s[696]), .cout(c[696]), .a(c[560]), .b(c[561]), .c(c[562]));
FA fa_3_21 (.sum(s[697]), .cout(c[697]), .a(s[563]), .b(s[564]), .c(s[565]));
FA fa_3_22 (.sum(s[698]), .cout(c[698]), .a(c[563]), .b(c[564]), .c(c[565]));
FA fa_3_23 (.sum(s[699]), .cout(c[699]), .a(s[566]), .b(s[567]), .c(s[568]));
FA fa_3_24 (.sum(s[700]), .cout(c[700]), .a(c[566]), .b(c[567]), .c(c[568]));
FA fa_3_25 (.sum(s[701]), .cout(c[701]), .a(s[569]), .b(s[570]), .c(s[571]));
FA fa_3_26 (.sum(s[702]), .cout(c[702]), .a(c[569]), .b(c[570]), .c(c[571]));
FA fa_3_27 (.sum(s[703]), .cout(c[703]), .a(s[572]), .b(s[573]), .c(s[574]));
FA fa_3_28 (.sum(s[704]), .cout(c[704]), .a(c[572]), .b(c[573]), .c(c[574]));
FA fa_3_29 (.sum(s[705]), .cout(c[705]), .a(c[575]), .b(s[576]), .c(s[577]));
FA fa_3_30 (.sum(s[706]), .cout(c[706]), .a(s[578]), .b(s[388]), .c(s[389]));
FA fa_3_31 (.sum(s[707]), .cout(c[707]), .a(c[576]), .b(c[577]), .c(c[578]));
FA fa_3_32 (.sum(s[708]), .cout(c[708]), .a(s[579]), .b(s[580]), .c(s[581]));
FA fa_3_33 (.sum(s[709]), .cout(c[709]), .a(c[579]), .b(c[580]), .c(c[581]));
FA fa_3_34 (.sum(s[710]), .cout(c[710]), .a(c[582]), .b(s[583]), .c(s[584]));
FA fa_3_35 (.sum(s[711]), .cout(c[711]), .a(c[583]), .b(c[584]), .c(c[585]));
FA fa_3_36 (.sum(s[712]), .cout(c[712]), .a(c[586]), .b(s[587]), .c(s[588]));
FA fa_3_37 (.sum(s[713]), .cout(c[713]), .a(s[589]), .b(s[590]), .c(p[27][1]));
FA fa_3_38 (.sum(s[714]), .cout(c[714]), .a(c[587]), .b(c[588]), .c(c[589]));
FA fa_3_39 (.sum(s[715]), .cout(c[715]), .a(c[590]), .b(s[591]), .c(s[592]));
FA fa_3_40 (.sum(s[716]), .cout(c[716]), .a(s[593]), .b(s[594]), .c(s[144]));
FA fa_3_41 (.sum(s[717]), .cout(c[717]), .a(c[591]), .b(c[592]), .c(c[593]));
FA fa_3_42 (.sum(s[718]), .cout(c[718]), .a(c[594]), .b(s[595]), .c(s[596]));
FA fa_3_43 (.sum(s[719]), .cout(c[719]), .a(s[597]), .b(s[598]), .c(s[419]));
FA fa_3_44 (.sum(s[720]), .cout(c[720]), .a(c[595]), .b(c[596]), .c(c[597]));
FA fa_3_45 (.sum(s[721]), .cout(c[721]), .a(c[598]), .b(s[599]), .c(s[600]));
FA fa_3_46 (.sum(s[722]), .cout(c[722]), .a(s[601]), .b(s[602]), .c(s[603]));
FA fa_3_47 (.sum(s[723]), .cout(c[723]), .a(c[599]), .b(c[600]), .c(c[601]));
FA fa_3_48 (.sum(s[724]), .cout(c[724]), .a(c[602]), .b(c[603]), .c(s[604]));
FA fa_3_49 (.sum(s[725]), .cout(c[725]), .a(s[605]), .b(s[606]), .c(s[607]));
FA fa_3_50 (.sum(s[726]), .cout(c[726]), .a(c[604]), .b(c[605]), .c(c[606]));
FA fa_3_51 (.sum(s[727]), .cout(c[727]), .a(c[607]), .b(s[608]), .c(s[609]));
FA fa_3_52 (.sum(s[728]), .cout(c[728]), .a(s[610]), .b(s[611]), .c(s[612]));
FA fa_3_53 (.sum(s[729]), .cout(c[729]), .a(c[608]), .b(c[609]), .c(c[610]));
FA fa_3_54 (.sum(s[730]), .cout(c[730]), .a(c[611]), .b(c[612]), .c(s[613]));
FA fa_3_55 (.sum(s[731]), .cout(c[731]), .a(s[614]), .b(s[615]), .c(s[616]));
FA fa_3_56 (.sum(s[732]), .cout(c[732]), .a(c[613]), .b(c[614]), .c(c[615]));
FA fa_3_57 (.sum(s[733]), .cout(c[733]), .a(c[616]), .b(s[617]), .c(s[618]));
FA fa_3_58 (.sum(s[734]), .cout(c[734]), .a(s[619]), .b(s[620]), .c(s[452]));
FA fa_3_59 (.sum(s[735]), .cout(c[735]), .a(c[617]), .b(c[618]), .c(c[619]));
FA fa_3_60 (.sum(s[736]), .cout(c[736]), .a(c[620]), .b(s[621]), .c(s[622]));
FA fa_3_61 (.sum(s[737]), .cout(c[737]), .a(c[621]), .b(c[622]), .c(c[623]));
FA fa_3_62 (.sum(s[738]), .cout(c[738]), .a(c[624]), .b(s[625]), .c(s[626]));
FA fa_3_63 (.sum(s[739]), .cout(c[739]), .a(s[627]), .b(s[628]), .c(p[31][6]));
FA fa_3_64 (.sum(s[740]), .cout(c[740]), .a(c[625]), .b(c[626]), .c(c[627]));
FA fa_3_65 (.sum(s[741]), .cout(c[741]), .a(c[628]), .b(s[629]), .c(s[630]));
FA fa_3_66 (.sum(s[742]), .cout(c[742]), .a(s[631]), .b(s[632]), .c(p[31][7]));
FA fa_3_67 (.sum(s[743]), .cout(c[743]), .a(c[629]), .b(c[630]), .c(c[631]));
FA fa_3_68 (.sum(s[744]), .cout(c[744]), .a(c[632]), .b(s[633]), .c(s[634]));
FA fa_3_69 (.sum(s[745]), .cout(c[745]), .a(s[635]), .b(s[474]), .c(s[235]));
FA fa_3_70 (.sum(s[746]), .cout(c[746]), .a(c[633]), .b(c[634]), .c(c[635]));
FA fa_3_71 (.sum(s[747]), .cout(c[747]), .a(s[636]), .b(s[637]), .c(s[638]));
FA fa_3_72 (.sum(s[748]), .cout(c[748]), .a(c[636]), .b(c[637]), .c(c[638]));
FA fa_3_73 (.sum(s[749]), .cout(c[749]), .a(c[639]), .b(s[640]), .c(s[641]));
FA fa_3_74 (.sum(s[750]), .cout(c[750]), .a(c[640]), .b(c[641]), .c(c[642]));
FA fa_3_75 (.sum(s[751]), .cout(c[751]), .a(s[643]), .b(s[644]), .c(s[645]));
FA fa_3_76 (.sum(s[752]), .cout(c[752]), .a(c[643]), .b(c[644]), .c(c[645]));
FA fa_3_77 (.sum(s[753]), .cout(c[753]), .a(s[646]), .b(s[647]), .c(s[648]));
FA fa_3_78 (.sum(s[754]), .cout(c[754]), .a(c[646]), .b(c[647]), .c(c[648]));
FA fa_3_79 (.sum(s[755]), .cout(c[755]), .a(s[649]), .b(s[650]), .c(s[651]));
FA fa_3_80 (.sum(s[756]), .cout(c[756]), .a(c[649]), .b(c[650]), .c(c[651]));
FA fa_3_81 (.sum(s[757]), .cout(c[757]), .a(s[652]), .b(s[653]), .c(s[500]));
FA fa_3_82 (.sum(s[758]), .cout(c[758]), .a(c[652]), .b(c[653]), .c(s[654]));
FA fa_3_83 (.sum(s[759]), .cout(c[759]), .a(c[654]), .b(c[655]), .c(c[656]));
FA fa_3_84 (.sum(s[760]), .cout(c[760]), .a(s[657]), .b(s[658]), .c(s[659]));
FA fa_3_85 (.sum(s[761]), .cout(c[761]), .a(c[657]), .b(c[658]), .c(c[659]));
FA fa_3_86 (.sum(s[762]), .cout(c[762]), .a(s[660]), .b(s[661]), .c(s[289]));
FA fa_3_87 (.sum(s[763]), .cout(c[763]), .a(c[660]), .b(c[661]), .c(s[662]));
FA fa_3_88 (.sum(s[764]), .cout(c[764]), .a(s[663]), .b(p[30][19]), .c(p[31][18]));
FA fa_3_89 (.sum(s[765]), .cout(c[765]), .a(c[662]), .b(c[663]), .c(s[664]));
FA fa_3_90 (.sum(s[766]), .cout(c[766]), .a(c[664]), .b(c[665]), .c(s[666]));
FA fa_3_91 (.sum(s[767]), .cout(c[767]), .a(c[666]), .b(c[667]), .c(s[668]));
FA fa_3_92 (.sum(s[768]), .cout(c[768]), .a(c[668]), .b(s[669]), .c(s[670]));
FA fa_3_93 (.sum(s[769]), .cout(c[769]), .a(c[669]), .b(c[670]), .c(s[671]));
FA fa_3_94 (.sum(s[770]), .cout(c[770]), .a(c[671]), .b(s[672]), .c(s[528]));
FA fa_3_95 (.sum(s[771]), .cout(c[771]), .a(c[672]), .b(s[673]), .c(s[314]));
FA fa_3_96 (.sum(s[772]), .cout(c[772]), .a(c[674]), .b(s[675]), .c(p[31][27]));
FA fa_3_97 (.sum(s[773]), .cout(c[773]), .a(c[675]), .b(c[531]), .c(s[532]));
HA ha_4_1 (.sum(s[774]), .cout(c[774]), .a(c[678]), .b(s[679]));
HA ha_4_2 (.sum(s[775]), .cout(c[775]), .a(c[679]), .b(s[680]));
HA ha_4_3 (.sum(s[776]), .cout(c[776]), .a(c[680]), .b(s[681]));
FA fa_4_4 (.sum(s[777]), .cout(c[777]), .a(c[681]), .b(s[682]), .c(s[332]));
FA fa_4_5 (.sum(s[778]), .cout(c[778]), .a(c[682]), .b(s[683]), .c(s[335]));
FA fa_4_6 (.sum(s[779]), .cout(c[779]), .a(c[683]), .b(s[684]), .c(p[13][0]));
FA fa_4_7 (.sum(s[780]), .cout(c[780]), .a(c[684]), .b(s[685]), .c(s[547]));
FA fa_4_8 (.sum(s[781]), .cout(c[781]), .a(c[685]), .b(s[686]), .c(s[687]));
FA fa_4_9 (.sum(s[782]), .cout(c[782]), .a(c[686]), .b(c[687]), .c(s[688]));
FA fa_4_10 (.sum(s[783]), .cout(c[783]), .a(c[688]), .b(s[689]), .c(s[553]));
FA fa_4_11 (.sum(s[784]), .cout(c[784]), .a(c[689]), .b(s[690]), .c(s[691]));
FA fa_4_12 (.sum(s[785]), .cout(c[785]), .a(c[690]), .b(c[691]), .c(s[692]));
FA fa_4_13 (.sum(s[786]), .cout(c[786]), .a(c[692]), .b(c[693]), .c(s[694]));
FA fa_4_14 (.sum(s[787]), .cout(c[787]), .a(c[694]), .b(c[695]), .c(s[696]));
FA fa_4_15 (.sum(s[788]), .cout(c[788]), .a(c[696]), .b(c[697]), .c(s[698]));
FA fa_4_16 (.sum(s[789]), .cout(c[789]), .a(s[699]), .b(s[373]), .c(p[22][0]));
FA fa_4_17 (.sum(s[790]), .cout(c[790]), .a(c[698]), .b(c[699]), .c(s[700]));
FA fa_4_18 (.sum(s[791]), .cout(c[791]), .a(c[700]), .b(c[701]), .c(s[702]));
FA fa_4_19 (.sum(s[792]), .cout(c[792]), .a(c[702]), .b(c[703]), .c(s[704]));
FA fa_4_20 (.sum(s[793]), .cout(c[793]), .a(c[704]), .b(c[705]), .c(c[706]));
FA fa_4_21 (.sum(s[794]), .cout(c[794]), .a(s[707]), .b(s[708]), .c(s[582]));
FA fa_4_22 (.sum(s[795]), .cout(c[795]), .a(c[707]), .b(c[708]), .c(s[709]));
FA fa_4_23 (.sum(s[796]), .cout(c[796]), .a(s[710]), .b(s[585]), .c(s[586]));
FA fa_4_24 (.sum(s[797]), .cout(c[797]), .a(c[709]), .b(c[710]), .c(s[711]));
FA fa_4_25 (.sum(s[798]), .cout(c[798]), .a(s[712]), .b(s[713]), .c(p[28][0]));
FA fa_4_26 (.sum(s[799]), .cout(c[799]), .a(c[711]), .b(c[712]), .c(c[713]));
FA fa_4_27 (.sum(s[800]), .cout(c[800]), .a(s[714]), .b(s[715]), .c(s[716]));
FA fa_4_28 (.sum(s[801]), .cout(c[801]), .a(c[714]), .b(c[715]), .c(c[716]));
FA fa_4_29 (.sum(s[802]), .cout(c[802]), .a(s[717]), .b(s[718]), .c(s[719]));
FA fa_4_30 (.sum(s[803]), .cout(c[803]), .a(c[717]), .b(c[718]), .c(c[719]));
FA fa_4_31 (.sum(s[804]), .cout(c[804]), .a(s[720]), .b(s[721]), .c(s[722]));
FA fa_4_32 (.sum(s[805]), .cout(c[805]), .a(c[720]), .b(c[721]), .c(c[722]));
FA fa_4_33 (.sum(s[806]), .cout(c[806]), .a(s[723]), .b(s[724]), .c(s[725]));
FA fa_4_34 (.sum(s[807]), .cout(c[807]), .a(c[723]), .b(c[724]), .c(c[725]));
FA fa_4_35 (.sum(s[808]), .cout(c[808]), .a(s[726]), .b(s[727]), .c(s[728]));
FA fa_4_36 (.sum(s[809]), .cout(c[809]), .a(c[726]), .b(c[727]), .c(c[728]));
FA fa_4_37 (.sum(s[810]), .cout(c[810]), .a(s[729]), .b(s[730]), .c(s[731]));
FA fa_4_38 (.sum(s[811]), .cout(c[811]), .a(c[729]), .b(c[730]), .c(c[731]));
FA fa_4_39 (.sum(s[812]), .cout(c[812]), .a(s[732]), .b(s[733]), .c(s[734]));
FA fa_4_40 (.sum(s[813]), .cout(c[813]), .a(c[732]), .b(c[733]), .c(c[734]));
FA fa_4_41 (.sum(s[814]), .cout(c[814]), .a(s[735]), .b(s[736]), .c(s[623]));
FA fa_4_42 (.sum(s[815]), .cout(c[815]), .a(c[735]), .b(c[736]), .c(s[737]));
FA fa_4_43 (.sum(s[816]), .cout(c[816]), .a(c[737]), .b(c[738]), .c(c[739]));
FA fa_4_44 (.sum(s[817]), .cout(c[817]), .a(s[740]), .b(s[741]), .c(s[742]));
FA fa_4_45 (.sum(s[818]), .cout(c[818]), .a(c[740]), .b(c[741]), .c(c[742]));
FA fa_4_46 (.sum(s[819]), .cout(c[819]), .a(s[743]), .b(s[744]), .c(s[745]));
FA fa_4_47 (.sum(s[820]), .cout(c[820]), .a(c[743]), .b(c[744]), .c(c[745]));
FA fa_4_48 (.sum(s[821]), .cout(c[821]), .a(s[746]), .b(s[747]), .c(s[639]));
FA fa_4_49 (.sum(s[822]), .cout(c[822]), .a(c[746]), .b(c[747]), .c(s[748]));
FA fa_4_50 (.sum(s[823]), .cout(c[823]), .a(s[749]), .b(s[642]), .c(s[484]));
FA fa_4_51 (.sum(s[824]), .cout(c[824]), .a(c[748]), .b(c[749]), .c(s[750]));
FA fa_4_52 (.sum(s[825]), .cout(c[825]), .a(s[751]), .b(s[255]), .c(s[256]));
FA fa_4_53 (.sum(s[826]), .cout(c[826]), .a(c[750]), .b(c[751]), .c(s[752]));
FA fa_4_54 (.sum(s[827]), .cout(c[827]), .a(c[752]), .b(c[753]), .c(s[754]));
FA fa_4_55 (.sum(s[828]), .cout(c[828]), .a(c[754]), .b(c[755]), .c(s[756]));
FA fa_4_56 (.sum(s[829]), .cout(c[829]), .a(c[756]), .b(c[757]), .c(s[758]));
FA fa_4_57 (.sum(s[830]), .cout(c[830]), .a(c[758]), .b(s[759]), .c(s[760]));
FA fa_4_58 (.sum(s[831]), .cout(c[831]), .a(c[759]), .b(c[760]), .c(s[761]));
FA fa_4_59 (.sum(s[832]), .cout(c[832]), .a(c[761]), .b(c[762]), .c(s[763]));
FA fa_4_60 (.sum(s[833]), .cout(c[833]), .a(c[763]), .b(c[764]), .c(s[765]));
FA fa_4_61 (.sum(s[834]), .cout(c[834]), .a(c[765]), .b(s[766]), .c(s[667]));
FA fa_4_62 (.sum(s[835]), .cout(c[835]), .a(c[766]), .b(s[767]), .c(s[521]));
FA fa_4_63 (.sum(s[836]), .cout(c[836]), .a(c[768]), .b(s[769]), .c(s[526]));
FA fa_4_64 (.sum(s[837]), .cout(c[837]), .a(c[769]), .b(s[770]), .c(p[31][24]));
FA fa_4_65 (.sum(s[838]), .cout(c[838]), .a(c[770]), .b(s[771]), .c(p[31][25]));
FA fa_4_66 (.sum(s[839]), .cout(c[839]), .a(c[771]), .b(c[673]), .c(s[674]));
HA ha_5_1 (.sum(s[840]), .cout(c[840]), .a(c[776]), .b(s[777]));
HA ha_5_2 (.sum(s[841]), .cout(c[841]), .a(c[777]), .b(s[778]));
HA ha_5_3 (.sum(s[842]), .cout(c[842]), .a(c[778]), .b(s[779]));
HA ha_5_4 (.sum(s[843]), .cout(c[843]), .a(c[779]), .b(s[780]));
HA ha_5_5 (.sum(s[844]), .cout(c[844]), .a(c[780]), .b(s[781]));
FA fa_5_6 (.sum(s[845]), .cout(c[845]), .a(c[781]), .b(s[782]), .c(s[551]));
FA fa_5_7 (.sum(s[846]), .cout(c[846]), .a(c[782]), .b(s[783]), .c(s[554]));
FA fa_5_8 (.sum(s[847]), .cout(c[847]), .a(c[783]), .b(s[784]), .c(p[18][0]));
FA fa_5_9 (.sum(s[848]), .cout(c[848]), .a(c[784]), .b(s[785]), .c(s[693]));
FA fa_5_10 (.sum(s[849]), .cout(c[849]), .a(c[785]), .b(s[786]), .c(s[695]));
FA fa_5_11 (.sum(s[850]), .cout(c[850]), .a(c[786]), .b(s[787]), .c(s[697]));
FA fa_5_12 (.sum(s[851]), .cout(c[851]), .a(c[787]), .b(s[788]), .c(s[789]));
FA fa_5_13 (.sum(s[852]), .cout(c[852]), .a(c[788]), .b(c[789]), .c(s[790]));
FA fa_5_14 (.sum(s[853]), .cout(c[853]), .a(c[790]), .b(s[791]), .c(s[703]));
FA fa_5_15 (.sum(s[854]), .cout(c[854]), .a(c[791]), .b(s[792]), .c(s[705]));
FA fa_5_16 (.sum(s[855]), .cout(c[855]), .a(c[792]), .b(s[793]), .c(s[794]));
FA fa_5_17 (.sum(s[856]), .cout(c[856]), .a(c[793]), .b(c[794]), .c(s[795]));
FA fa_5_18 (.sum(s[857]), .cout(c[857]), .a(c[795]), .b(c[796]), .c(s[797]));
FA fa_5_19 (.sum(s[858]), .cout(c[858]), .a(c[797]), .b(c[798]), .c(s[799]));
FA fa_5_20 (.sum(s[859]), .cout(c[859]), .a(c[799]), .b(c[800]), .c(s[801]));
FA fa_5_21 (.sum(s[860]), .cout(c[860]), .a(c[801]), .b(c[802]), .c(s[803]));
FA fa_5_22 (.sum(s[861]), .cout(c[861]), .a(c[803]), .b(c[804]), .c(s[805]));
FA fa_5_23 (.sum(s[862]), .cout(c[862]), .a(s[806]), .b(s[432]), .c(s[433]));
FA fa_5_24 (.sum(s[863]), .cout(c[863]), .a(c[805]), .b(c[806]), .c(s[807]));
FA fa_5_25 (.sum(s[864]), .cout(c[864]), .a(c[807]), .b(c[808]), .c(s[809]));
FA fa_5_26 (.sum(s[865]), .cout(c[865]), .a(c[809]), .b(c[810]), .c(s[811]));
FA fa_5_27 (.sum(s[866]), .cout(c[866]), .a(c[811]), .b(c[812]), .c(s[813]));
FA fa_5_28 (.sum(s[867]), .cout(c[867]), .a(c[813]), .b(c[814]), .c(s[815]));
FA fa_5_29 (.sum(s[868]), .cout(c[868]), .a(c[815]), .b(s[816]), .c(s[817]));
FA fa_5_30 (.sum(s[869]), .cout(c[869]), .a(c[816]), .b(c[817]), .c(s[818]));
FA fa_5_31 (.sum(s[870]), .cout(c[870]), .a(c[818]), .b(c[819]), .c(s[820]));
FA fa_5_32 (.sum(s[871]), .cout(c[871]), .a(c[820]), .b(c[821]), .c(s[822]));
FA fa_5_33 (.sum(s[872]), .cout(c[872]), .a(c[822]), .b(c[823]), .c(s[824]));
FA fa_5_34 (.sum(s[873]), .cout(c[873]), .a(c[824]), .b(c[825]), .c(s[826]));
FA fa_5_35 (.sum(s[874]), .cout(c[874]), .a(c[826]), .b(s[827]), .c(s[755]));
FA fa_5_36 (.sum(s[875]), .cout(c[875]), .a(c[827]), .b(s[828]), .c(s[757]));
FA fa_5_37 (.sum(s[876]), .cout(c[876]), .a(c[828]), .b(s[829]), .c(s[655]));
FA fa_5_38 (.sum(s[877]), .cout(c[877]), .a(c[830]), .b(s[831]), .c(s[762]));
FA fa_5_39 (.sum(s[878]), .cout(c[878]), .a(c[831]), .b(s[832]), .c(s[764]));
FA fa_5_40 (.sum(s[879]), .cout(c[879]), .a(c[832]), .b(s[833]), .c(s[665]));
FA fa_5_41 (.sum(s[880]), .cout(c[880]), .a(c[833]), .b(s[834]), .c(s[301]));
FA fa_5_42 (.sum(s[881]), .cout(c[881]), .a(c[834]), .b(s[835]), .c(s[522]));
FA fa_5_43 (.sum(s[882]), .cout(c[882]), .a(c[835]), .b(c[767]), .c(s[768]));
HA ha_6_1 (.sum(s[883]), .cout(c[883]), .a(c[844]), .b(s[845]));
HA ha_6_2 (.sum(s[884]), .cout(c[884]), .a(c[845]), .b(s[846]));
HA ha_6_3 (.sum(s[885]), .cout(c[885]), .a(c[846]), .b(s[847]));
HA ha_6_4 (.sum(s[886]), .cout(c[886]), .a(c[847]), .b(s[848]));
HA ha_6_5 (.sum(s[887]), .cout(c[887]), .a(c[848]), .b(s[849]));
HA ha_6_6 (.sum(s[888]), .cout(c[888]), .a(c[849]), .b(s[850]));
HA ha_6_7 (.sum(s[889]), .cout(c[889]), .a(c[850]), .b(s[851]));
FA fa_6_8 (.sum(s[890]), .cout(c[890]), .a(c[851]), .b(s[852]), .c(s[701]));
FA fa_6_9 (.sum(s[891]), .cout(c[891]), .a(c[852]), .b(s[853]), .c(s[575]));
FA fa_6_10 (.sum(s[892]), .cout(c[892]), .a(c[853]), .b(s[854]), .c(s[706]));
FA fa_6_11 (.sum(s[893]), .cout(c[893]), .a(c[854]), .b(s[855]), .c(s[116]));
FA fa_6_12 (.sum(s[894]), .cout(c[894]), .a(c[855]), .b(s[856]), .c(s[796]));
FA fa_6_13 (.sum(s[895]), .cout(c[895]), .a(c[856]), .b(s[857]), .c(s[798]));
FA fa_6_14 (.sum(s[896]), .cout(c[896]), .a(c[857]), .b(s[858]), .c(s[800]));
FA fa_6_15 (.sum(s[897]), .cout(c[897]), .a(c[858]), .b(s[859]), .c(s[802]));
FA fa_6_16 (.sum(s[898]), .cout(c[898]), .a(c[859]), .b(s[860]), .c(s[804]));
FA fa_6_17 (.sum(s[899]), .cout(c[899]), .a(c[860]), .b(s[861]), .c(s[862]));
FA fa_6_18 (.sum(s[900]), .cout(c[900]), .a(c[861]), .b(c[862]), .c(s[863]));
FA fa_6_19 (.sum(s[901]), .cout(c[901]), .a(c[863]), .b(s[864]), .c(s[810]));
FA fa_6_20 (.sum(s[902]), .cout(c[902]), .a(c[864]), .b(s[865]), .c(s[812]));
FA fa_6_21 (.sum(s[903]), .cout(c[903]), .a(c[865]), .b(s[866]), .c(s[814]));
FA fa_6_22 (.sum(s[904]), .cout(c[904]), .a(c[866]), .b(s[867]), .c(s[738]));
FA fa_6_23 (.sum(s[905]), .cout(c[905]), .a(c[868]), .b(s[869]), .c(s[819]));
FA fa_6_24 (.sum(s[906]), .cout(c[906]), .a(c[869]), .b(s[870]), .c(s[821]));
FA fa_6_25 (.sum(s[907]), .cout(c[907]), .a(c[870]), .b(s[871]), .c(s[823]));
FA fa_6_26 (.sum(s[908]), .cout(c[908]), .a(c[871]), .b(s[872]), .c(s[825]));
FA fa_6_27 (.sum(s[909]), .cout(c[909]), .a(c[872]), .b(s[873]), .c(s[753]));
FA fa_6_28 (.sum(s[910]), .cout(c[910]), .a(c[873]), .b(s[874]), .c(p[31][13]));
FA fa_6_29 (.sum(s[911]), .cout(c[911]), .a(c[874]), .b(s[875]), .c(s[501]));
FA fa_6_30 (.sum(s[912]), .cout(c[912]), .a(c[875]), .b(s[876]), .c(s[656]));
FA fa_6_31 (.sum(s[913]), .cout(c[913]), .a(c[876]), .b(c[829]), .c(s[830]));
HA ha_7_1 (.sum(s[914]), .cout(c[914]), .a(c[889]), .b(s[890]));
HA ha_7_2 (.sum(s[915]), .cout(c[915]), .a(c[890]), .b(s[891]));
HA ha_7_3 (.sum(s[916]), .cout(c[916]), .a(c[891]), .b(s[892]));
HA ha_7_4 (.sum(s[917]), .cout(c[917]), .a(c[892]), .b(s[893]));
HA ha_7_5 (.sum(s[918]), .cout(c[918]), .a(c[893]), .b(s[894]));
HA ha_7_6 (.sum(s[919]), .cout(c[919]), .a(c[894]), .b(s[895]));
HA ha_7_7 (.sum(s[920]), .cout(c[920]), .a(c[895]), .b(s[896]));
HA ha_7_8 (.sum(s[921]), .cout(c[921]), .a(c[896]), .b(s[897]));
HA ha_7_9 (.sum(s[922]), .cout(c[922]), .a(c[897]), .b(s[898]));
HA ha_7_10 (.sum(s[923]), .cout(c[923]), .a(c[898]), .b(s[899]));
FA fa_7_11 (.sum(s[924]), .cout(c[924]), .a(c[899]), .b(s[900]), .c(s[808]));
FA fa_7_12 (.sum(s[925]), .cout(c[925]), .a(c[900]), .b(s[901]), .c(s[446]));
FA fa_7_13 (.sum(s[926]), .cout(c[926]), .a(c[901]), .b(s[902]), .c(p[31][4]));
FA fa_7_14 (.sum(s[927]), .cout(c[927]), .a(c[902]), .b(s[903]), .c(s[624]));
FA fa_7_15 (.sum(s[928]), .cout(c[928]), .a(c[903]), .b(s[904]), .c(s[739]));
FA fa_7_16 (.sum(s[929]), .cout(c[929]), .a(c[904]), .b(c[867]), .c(s[868]));

endmodule