module datamux(
    input logic[255:0] data_one,
    input logic[255:0] data_two,
    input logic[4:0] offset,
    input logic use_set_one,

    output logic[32:0] out
    );






endmodule
